
    `ifndef CIRC_SPEC_gb4
    `define CIRC_SPEC_gb4
    localparam integer NUM_CONSTS = 4;
    localparam integer NUM_VARS = 16;
    localparam integer NUM_OUTPUTS = 4;

    localparam integer NUM_INPUTS = NUM_CONSTS + NUM_VARS;
    localparam integer NUM_WEIGHTS = 2 ** NUM_VARS;
    localparam integer WEIGHT_MATRIX [NUM_OUTPUTS * NUM_WEIGHTS-1 : 0]   = {0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,0,1,2,3,1,2,3,4,0,1,2,3,1,2,3,4,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,1,2,3,4,2,3,4,5,1,2,3,4,2,3,4,5,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,2,3,4,5,3,4,5,6,2,3,4,5,3,4,5,6,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,3,4,5,6,4,5,6,7,3,4,5,6,4,5,6,7,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,5,6,7,8,6,7,8,9,5,6,7,8,6,7,8,9,7,8,9,10,8,9,10,11,7,8,9,10,8,9,10,11,9,10,11,12,10,11,12,13,9,10,11,12,10,11,12,13,11,12,13,14,12,13,14,15,11,12,13,14,12,13,14,15,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,4,5,6,7,5,6,7,8,4,5,6,7,5,6,7,8,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,6,7,8,9,7,8,9,10,6,7,8,9,7,8,9,10,8,9,10,11,9,10,11,12,8,9,10,11,9,10,11,12,10,11,12,13,11,12,13,14,10,11,12,13,11,12,13,14,12,13,14,15,13,14,15,16,12,13,14,15,13,14,15,16,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,0,0,1,1,2,2,3,3,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,1,1,2,2,3,3,4,4,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,2,2,3,3,4,4,5,5,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,3,3,4,4,5,5,6,6,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,4,4,5,5,6,6,7,7,5,5,6,6,7,7,8,8,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,6,6,7,7,8,8,9,9,7,7,8,8,9,9,10,10,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,8,8,9,9,10,10,11,11,9,9,10,10,11,11,12,12,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,10,10,11,11,12,12,13,13,11,11,12,12,13,13,14,14,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,12,12,13,13,14,14,15,15,13,13,14,14,15,15,16,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16};
    `endif
    