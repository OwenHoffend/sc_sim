`define HMT_IMPLEMENTATION
`ifdef HMT_IMPLEMENTATION
module mux_1(
	input s, x, y,
	output logic z
);
	assign z = s ? y : x;
endmodule

module gb3_linear(
	input  x1, x2, x3, c0, c1,
	output logic z
);
	logic a1;
	mux_1 m1(c0, x1, x3, a1);
	mux_1 m2(c1, a1, x2, z);
endmodule

module gb3(
    input x11, x12, x13,
          x21, x22, x23,
          x31, x32, x33,
          c0, c1, c2, c3,
	output logic z
);
	logic a1, a2, a3;
    gb3_linear gb3_1(x11, x12, x13, c0, c1, a1);
    gb3_linear gb3_2(x21, x22, x23, c0, c1, a2);
    gb3_linear gb3_3(x31, x32, x33, c0, c1, a3);
	gb3_linear gb3_4(a1, a2, a3, c2, c3, z);
endmodule
`endif

module gb4(
    input [19:0] x,
    output logic [3:0] z
);

`ifdef HMT_IMPLEMENTATION

logic x11, x12, x13, x14,
    x21, x22, x23, x24,
    x31, x32, x33, x34,
    x41, x42, x43, x44,
    c0, c1, c2, c3;

assign x11 = x[19];
assign x12 = x[18];
assign x13 = x[17];
assign x14 = x[16];
assign x21 = x[15];
assign x22 = x[14];
assign x23 = x[13];
assign x24 = x[12];
assign x31 = x[11];
assign x32 = x[10];
assign x33 = x[9];
assign x34 = x[8];
assign x41 = x[7];
assign x42 = x[6];
assign x43 = x[5];
assign x44 = x[4];
assign c0 = x[3];
assign c1 = x[2];
assign c2 = x[1];
assign c3 = x[0];

    gb3 gb3_1( //ul (x11)
        x11, x12, x13,
        x21, x22, x23,
        x31, x32, x33,
        c0, c1, c2, c3,
        z[0]
    );
    gb3 gb3_2( //ur (x12)
        x12, x13, x14,
        x22, x23, x24,
        x32, x33, x34,
        c0, c1, c2, c3,
        z[1]
    );
    gb3 gb3_3( //ll (x21)
        x21, x22, x23,
        x31, x32, x33,
        x41, x42, x43,
        c0, c1, c2, c3,
        z[2]
    );
    gb3 gb3_4( //lr (x22)
        x22, x23, x24,
        x32, x33, x34,
        x42, x43, x44,
        c0, c1, c2, c3,
        z[3]
    );
`else
always_comb begin 
	 z = 4'b0000;
	if(x==?20'b111?111?111?????????) z |= 4'b1000; 
	if(x==?20'b?111?111?111????????) z |= 4'b0100; 
	if(x==?20'b????111?111?111?????) z |= 4'b0010; 
	if(x==?20'b?????111?111?111????) z |= 4'b0001; 
	if(x==?20'b111?????111????????1) z |= 4'b1000; 
	if(x==?20'b?111?????111???????1) z |= 4'b0100; 
	if(x==?20'b????111?????111????1) z |= 4'b0010; 
	if(x==?20'b?????111?????111???1) z |= 4'b0001; 
	if(x==?20'b111?111???????????1?) z |= 4'b1000; 
	if(x==?20'b?111?111??????????1?) z |= 4'b0100; 
	if(x==?20'b????????111?111???1?) z |= 4'b0010; 
	if(x==?20'b?????????111?111??1?) z |= 4'b0001; 
	if(x==?20'b11??11??11??????1???) z |= 4'b1000; 
	if(x==?20'b??11??11??11????1???) z |= 4'b0100; 
	if(x==?20'b????11??11??11??1???) z |= 4'b0010; 
	if(x==?20'b??????11??11??111???) z |= 4'b0001; 
	if(x==?20'b1?1?1?1?1?1??????1??) z |= 4'b1000; 
	if(x==?20'b?1?1?1?1?1?1?????1??) z |= 4'b0100; 
	if(x==?20'b????1?1?1?1?1?1??1??) z |= 4'b0010; 
	if(x==?20'b?????1?1?1?1?1?1?1??) z |= 4'b0001; 
	if(x==?20'b?11?11??11??????1???) z |= 4'b1000; 
	if(x==?20'b?11???11??11????1???) z |= 4'b0100; 
	if(x==?20'b????11??11???11?1???) z |= 4'b0010; 
	if(x==?20'b??????11??11?11?1???) z |= 4'b0001; 
	if(x==?20'b11??11???11?????1???) z |= 4'b1000; 
	if(x==?20'b11???11?11??????1???) z |= 4'b1000; 
	if(x==?20'b??11?11???11????1???) z |= 4'b0100; 
	if(x==?20'b??11??11?11?????1???) z |= 4'b0100; 
	if(x==?20'b????11???11?11??1???) z |= 4'b0010; 
	if(x==?20'b?????11?11??11??1???) z |= 4'b0010; 
	if(x==?20'b?????11???11??111???) z |= 4'b0001; 
	if(x==?20'b??????11?11???111???) z |= 4'b0001; 
	if(x==?20'b?11?11???11?????1???) z |= 4'b1000; 
	if(x==?20'b?11??11?11??????1???) z |= 4'b1000; 
	if(x==?20'b?11??11???11????1???) z |= 4'b0100; 
	if(x==?20'b?11???11?11?????1???) z |= 4'b0100; 
	if(x==?20'b????11???11??11?1???) z |= 4'b0010; 
	if(x==?20'b?????11?11???11?1???) z |= 4'b0010; 
	if(x==?20'b?????11???11?11?1???) z |= 4'b0001; 
	if(x==?20'b??????11?11??11?1???) z |= 4'b0001; 
	if(x==?20'b11???11??11?????1???) z |= 4'b1000; 
	if(x==?20'b??11?11??11?????1???) z |= 4'b0100; 
	if(x==?20'b?????11??11?11??1???) z |= 4'b0010; 
	if(x==?20'b?????11??11???111???) z |= 4'b0001; 
	if(x==?20'b????111?111???????1?) z |= 4'b1010; 
	if(x==?20'b?????111?111??????1?) z |= 4'b0101; 
	if(x==?20'b?11??11??11?????1???) z |= 4'b1100; 
	if(x==?20'b?????11??11??11?1???) z |= 4'b0011; 
	if(x==?20'b11??????11??????1??1) z |= 4'b1000; 
	if(x==?20'b??11??????11????1??1) z |= 4'b0100; 
	if(x==?20'b????11??????11??1??1) z |= 4'b0010; 
	if(x==?20'b??????11??????111??1) z |= 4'b0001; 
	if(x==?20'b1?1??1??1?1??????1??) z |= 4'b1000; 
	if(x==?20'b1?1?1?1??1???????1??) z |= 4'b1000; 
	if(x==?20'b?1?1??1??1?1?????1??) z |= 4'b0100; 
	if(x==?20'b?1?1?1?1??1??????1??) z |= 4'b0100; 
	if(x==?20'b?????1??1?1?1?1??1??) z |= 4'b0010; 
	if(x==?20'b????1?1??1??1?1??1??) z |= 4'b0010; 
	if(x==?20'b??????1??1?1?1?1?1??) z |= 4'b0001; 
	if(x==?20'b?????1?1??1??1?1?1??) z |= 4'b0001; 
	if(x==?20'b11??11??????????1?1?) z |= 4'b1000; 
	if(x==?20'b??11??11????????1?1?) z |= 4'b0100; 
	if(x==?20'b????????11??11??1?1?) z |= 4'b0010; 
	if(x==?20'b??????????11??111?1?) z |= 4'b0001; 
	if(x==?20'b1?1?????1?1??????1?1) z |= 4'b1000; 
	if(x==?20'b?1?1?????1?1?????1?1) z |= 4'b0100; 
	if(x==?20'b????1?1?????1?1??1?1) z |= 4'b0010; 
	if(x==?20'b?????1?1?????1?1?1?1) z |= 4'b0001; 
	if(x==?20'b1?1?1?1??????????11?) z |= 4'b1000; 
	if(x==?20'b?1?1?1?1?????????11?) z |= 4'b0100; 
	if(x==?20'b????????1?1?1?1??11?) z |= 4'b0010; 
	if(x==?20'b?????????1?1?1?1?11?) z |= 4'b0001; 
	if(x==?20'b?1??1?1?1?1??????1??) z |= 4'b1000; 
	if(x==?20'b??1??1?1?1?1?????1??) z |= 4'b0100; 
	if(x==?20'b????1?1?1?1??1???1??) z |= 4'b0010; 
	if(x==?20'b?????1?1?1?1??1??1??) z |= 4'b0001; 
	if(x==?20'b?11?????11??????1??1) z |= 4'b1000; 
	if(x==?20'b?11???????11????1??1) z |= 4'b0100; 
	if(x==?20'b????11???????11?1??1) z |= 4'b0010; 
	if(x==?20'b??????11?????11?1??1) z |= 4'b0001; 
	if(x==?20'b?11?11??????????1?1?) z |= 4'b1000; 
	if(x==?20'b?11???11????????1?1?) z |= 4'b0100; 
	if(x==?20'b????????11???11?1?1?) z |= 4'b0010; 
	if(x==?20'b??????????11?11?1?1?) z |= 4'b0001; 
	if(x==?20'b11???????11?????1??1) z |= 4'b1000; 
	if(x==?20'b??11?????11?????1??1) z |= 4'b0100; 
	if(x==?20'b?????11?????11??1??1) z |= 4'b0010; 
	if(x==?20'b?????11???????111??1) z |= 4'b0001; 
	if(x==?20'b11???11?????????1?1?) z |= 4'b1000; 
	if(x==?20'b??11?11?????????1?1?) z |= 4'b0100; 
	if(x==?20'b?????????11?11??1?1?) z |= 4'b0010; 
	if(x==?20'b?????????11???111?1?) z |= 4'b0001; 
	if(x==?20'b111???????????????11) z |= 4'b1000; 
	if(x==?20'b?111??????????????11) z |= 4'b0100; 
	if(x==?20'b????????????111???11) z |= 4'b0010; 
	if(x==?20'b?????????????111??11) z |= 4'b0001; 
	if(x==?20'b????11??11??????1?1?) z |= 4'b1010; 
	if(x==?20'b??????11??11????1?1?) z |= 4'b0101; 
	if(x==?20'b?11??????11?????1??1) z |= 4'b1100; 
	if(x==?20'b?????11??????11?1??1) z |= 4'b0011; 
	if(x==?20'b?11??11?????????1?1?) z |= 4'b1100; 
	if(x==?20'b?????????11??11?1?1?) z |= 4'b0011; 
	if(x==?20'b????1?1?1?1??????11?) z |= 4'b1010; 
	if(x==?20'b?????1?1?1?1?????11?) z |= 4'b0101; 
	if(x==?20'b????11???11?????1?1?) z |= 4'b1010; 
	if(x==?20'b?????11?11??????1?1?) z |= 4'b1010; 
	if(x==?20'b?????11???11????1?1?) z |= 4'b0101; 
	if(x==?20'b??????11?11?????1?1?) z |= 4'b0101; 
	if(x==?20'b????????111???????11) z |= 4'b1000; 
	if(x==?20'b?????????111??????11) z |= 4'b0100; 
	if(x==?20'b????111???????????11) z |= 4'b0010; 
	if(x==?20'b?????111??????????11) z |= 4'b0001; 
	if(x==?20'b1?1??1???1???????1??) z |= 4'b1000; 
	if(x==?20'b?1?1??1???1??????1??) z |= 4'b0100; 
	if(x==?20'b?????1???1??1?1??1??) z |= 4'b0010; 
	if(x==?20'b??????1???1??1?1?1??) z |= 4'b0001; 
	if(x==?20'b1?1??????1???????1?1) z |= 4'b1000; 
	if(x==?20'b?1?1??????1??????1?1) z |= 4'b0100; 
	if(x==?20'b?????1??????1?1??1?1) z |= 4'b0010; 
	if(x==?20'b??????1??????1?1?1?1) z |= 4'b0001; 
	if(x==?20'b11??????????????1?11) z |= 4'b1000; 
	if(x==?20'b??11????????????1?11) z |= 4'b0100; 
	if(x==?20'b????????????11??1?11) z |= 4'b0010; 
	if(x==?20'b??????????????111?11) z |= 4'b0001; 
	if(x==?20'b1?1??1???????????11?) z |= 4'b1000; 
	if(x==?20'b?1?1??1??????????11?) z |= 4'b0100; 
	if(x==?20'b?????????1??1?1??11?) z |= 4'b0010; 
	if(x==?20'b??????????1??1?1?11?) z |= 4'b0001; 
	if(x==?20'b1?1??????????????111) z |= 4'b1000; 
	if(x==?20'b?1?1?????????????111) z |= 4'b0100; 
	if(x==?20'b????????????1?1??111) z |= 4'b0010; 
	if(x==?20'b?????????????1?1?111) z |= 4'b0001; 
	if(x==?20'b?1???1??1?1??????1??) z |= 4'b1000; 
	if(x==?20'b?1??1?1??1???????1??) z |= 4'b1000; 
	if(x==?20'b??1???1??1?1?????1??) z |= 4'b0100; 
	if(x==?20'b??1??1?1??1??????1??) z |= 4'b0100; 
	if(x==?20'b?????1??1?1??1???1??) z |= 4'b0010; 
	if(x==?20'b????1?1??1???1???1??) z |= 4'b0010; 
	if(x==?20'b??????1??1?1??1??1??) z |= 4'b0001; 
	if(x==?20'b?????1?1??1???1??1??) z |= 4'b0001; 
	if(x==?20'b?1??????1?1??????1?1) z |= 4'b1000; 
	if(x==?20'b??1??????1?1?????1?1) z |= 4'b0100; 
	if(x==?20'b????1?1??????1???1?1) z |= 4'b0010; 
	if(x==?20'b?????1?1??????1??1?1) z |= 4'b0001; 
	if(x==?20'b?1??1?1??????????11?) z |= 4'b1000; 
	if(x==?20'b??1??1?1?????????11?) z |= 4'b0100; 
	if(x==?20'b????????1?1??1???11?) z |= 4'b0010; 
	if(x==?20'b?????????1?1??1??11?) z |= 4'b0001; 
	if(x==?20'b1???1???1???????11??) z |= 4'b1000; 
	if(x==?20'b???1???1???1????11??) z |= 4'b0100; 
	if(x==?20'b????1???1???1???11??) z |= 4'b0010; 
	if(x==?20'b???????1???1???111??) z |= 4'b0001; 
	if(x==?20'b????????11??????1?11) z |= 4'b1000; 
	if(x==?20'b??????????11????1?11) z |= 4'b0100; 
	if(x==?20'b????11??????????1?11) z |= 4'b0010; 
	if(x==?20'b??????11????????1?11) z |= 4'b0001; 
	if(x==?20'b??1?1???1???????11??) z |= 4'b1000; 
	if(x==?20'b?1??1???1???????11??) z |= 4'b1000; 
	if(x==?20'b??1????1???1????11??) z |= 4'b0100; 
	if(x==?20'b?1?????1???1????11??) z |= 4'b0100; 
	if(x==?20'b????1???1?????1?11??) z |= 4'b0010; 
	if(x==?20'b????1???1????1??11??) z |= 4'b0010; 
	if(x==?20'b???????1???1??1?11??) z |= 4'b0001; 
	if(x==?20'b???????1???1?1??11??) z |= 4'b0001; 
	if(x==?20'b????????1?1??????111) z |= 4'b1000; 
	if(x==?20'b?????????1?1?????111) z |= 4'b0100; 
	if(x==?20'b????1?1??????????111) z |= 4'b0010; 
	if(x==?20'b?????1?1?????????111) z |= 4'b0001; 
	if(x==?20'b1???1?????1?????11??) z |= 4'b1000; 
	if(x==?20'b1???1????1??????11??) z |= 4'b1000; 
	if(x==?20'b1?????1?1???????11??) z |= 4'b1000; 
	if(x==?20'b1????1??1???????11??) z |= 4'b1000; 
	if(x==?20'b???1??1????1????11??) z |= 4'b0100; 
	if(x==?20'b???1?1?????1????11??) z |= 4'b0100; 
	if(x==?20'b???1???1??1?????11??) z |= 4'b0100; 
	if(x==?20'b???1???1?1??????11??) z |= 4'b0100; 
	if(x==?20'b????1?????1?1???11??) z |= 4'b0010; 
	if(x==?20'b????1????1??1???11??) z |= 4'b0010; 
	if(x==?20'b??????1?1???1???11??) z |= 4'b0010; 
	if(x==?20'b?????1??1???1???11??) z |= 4'b0010; 
	if(x==?20'b??????1????1???111??) z |= 4'b0001; 
	if(x==?20'b?????1?????1???111??) z |= 4'b0001; 
	if(x==?20'b???????1??1????111??) z |= 4'b0001; 
	if(x==?20'b???????1?1?????111??) z |= 4'b0001; 
	if(x==?20'b1???????1???????11?1) z |= 4'b1000; 
	if(x==?20'b???1???????1????11?1) z |= 4'b0100; 
	if(x==?20'b????1???????1???11?1) z |= 4'b0010; 
	if(x==?20'b???????1???????111?1) z |= 4'b0001; 
	if(x==?20'b1???1???????????111?) z |= 4'b1000; 
	if(x==?20'b???1???1????????111?) z |= 4'b0100; 
	if(x==?20'b????????1???1???111?) z |= 4'b0010; 
	if(x==?20'b???????????1???1111?) z |= 4'b0001; 
	if(x==?20'b?11?????????????1?11) z |= 4'b1100; 
	if(x==?20'b?????????????11?1?11) z |= 4'b0011; 
	if(x==?20'b??1?1?????1?????11??) z |= 4'b1000; 
	if(x==?20'b?1??1?????1?????11??) z |= 4'b1000; 
	if(x==?20'b??1?1????1??????11??) z |= 4'b1000; 
	if(x==?20'b?1??1????1??????11??) z |= 4'b1000; 
	if(x==?20'b??1???1?1???????11??) z |= 4'b1000; 
	if(x==?20'b?1????1?1???????11??) z |= 4'b1000; 
	if(x==?20'b??1??1??1???????11??) z |= 4'b1000; 
	if(x==?20'b?1???1??1???????11??) z |= 4'b1000; 
	if(x==?20'b??1???1????1????11??) z |= 4'b0100; 
	if(x==?20'b?1????1????1????11??) z |= 4'b0100; 
	if(x==?20'b??1??1?????1????11??) z |= 4'b0100; 
	if(x==?20'b?1???1?????1????11??) z |= 4'b0100; 
	if(x==?20'b??1????1??1?????11??) z |= 4'b0100; 
	if(x==?20'b?1?????1??1?????11??) z |= 4'b0100; 
	if(x==?20'b??1????1?1??????11??) z |= 4'b0100; 
	if(x==?20'b?1?????1?1??????11??) z |= 4'b0100; 
	if(x==?20'b????1?????1???1?11??) z |= 4'b0010; 
	if(x==?20'b????1????1????1?11??) z |= 4'b0010; 
	if(x==?20'b??????1?1?????1?11??) z |= 4'b0010; 
	if(x==?20'b?????1??1?????1?11??) z |= 4'b0010; 
	if(x==?20'b????1?????1??1??11??) z |= 4'b0010; 
	if(x==?20'b????1????1???1??11??) z |= 4'b0010; 
	if(x==?20'b??????1?1????1??11??) z |= 4'b0010; 
	if(x==?20'b?????1??1????1??11??) z |= 4'b0010; 
	if(x==?20'b??????1????1??1?11??) z |= 4'b0001; 
	if(x==?20'b?????1?????1??1?11??) z |= 4'b0001; 
	if(x==?20'b???????1??1???1?11??) z |= 4'b0001; 
	if(x==?20'b???????1?1????1?11??) z |= 4'b0001; 
	if(x==?20'b??????1????1?1??11??) z |= 4'b0001; 
	if(x==?20'b?????1?????1?1??11??) z |= 4'b0001; 
	if(x==?20'b???????1??1??1??11??) z |= 4'b0001; 
	if(x==?20'b???????1?1???1??11??) z |= 4'b0001; 
	if(x==?20'b??1?????1???????11?1) z |= 4'b1000; 
	if(x==?20'b?1??????1???????11?1) z |= 4'b1000; 
	if(x==?20'b??1????????1????11?1) z |= 4'b0100; 
	if(x==?20'b?1?????????1????11?1) z |= 4'b0100; 
	if(x==?20'b????1?????????1?11?1) z |= 4'b0010; 
	if(x==?20'b????1????????1??11?1) z |= 4'b0010; 
	if(x==?20'b???????1??????1?11?1) z |= 4'b0001; 
	if(x==?20'b???????1?????1??11?1) z |= 4'b0001; 
	if(x==?20'b??1?1???????????111?) z |= 4'b1000; 
	if(x==?20'b?1??1???????????111?) z |= 4'b1000; 
	if(x==?20'b??1????1????????111?) z |= 4'b0100; 
	if(x==?20'b?1?????1????????111?) z |= 4'b0100; 
	if(x==?20'b????????1?????1?111?) z |= 4'b0010; 
	if(x==?20'b????????1????1??111?) z |= 4'b0010; 
	if(x==?20'b???????????1??1?111?) z |= 4'b0001; 
	if(x==?20'b???????????1?1??111?) z |= 4'b0001; 
	if(x==?20'b1?????1???1?????11??) z |= 4'b1000; 
	if(x==?20'b1????1????1?????11??) z |= 4'b1000; 
	if(x==?20'b1?????1??1??????11??) z |= 4'b1000; 
	if(x==?20'b1????1???1??????11??) z |= 4'b1000; 
	if(x==?20'b???1??1???1?????11??) z |= 4'b0100; 
	if(x==?20'b???1?1????1?????11??) z |= 4'b0100; 
	if(x==?20'b???1??1??1??????11??) z |= 4'b0100; 
	if(x==?20'b???1?1???1??????11??) z |= 4'b0100; 
	if(x==?20'b??????1???1?1???11??) z |= 4'b0010; 
	if(x==?20'b?????1????1?1???11??) z |= 4'b0010; 
	if(x==?20'b??????1??1??1???11??) z |= 4'b0010; 
	if(x==?20'b?????1???1??1???11??) z |= 4'b0010; 
	if(x==?20'b??????1???1????111??) z |= 4'b0001; 
	if(x==?20'b?????1????1????111??) z |= 4'b0001; 
	if(x==?20'b??????1??1?????111??) z |= 4'b0001; 
	if(x==?20'b?????1???1?????111??) z |= 4'b0001; 
	if(x==?20'b????111????????????1) z |= 4'b1000; 
	if(x==?20'b?????111???????????1) z |= 4'b0100; 
	if(x==?20'b????????111????????1) z |= 4'b0010; 
	if(x==?20'b?????????111???????1) z |= 4'b0001; 
	if(x==?20'b1?????????1?????11?1) z |= 4'b1000; 
	if(x==?20'b1????????1??????11?1) z |= 4'b1000; 
	if(x==?20'b???1??????1?????11?1) z |= 4'b0100; 
	if(x==?20'b???1?????1??????11?1) z |= 4'b0100; 
	if(x==?20'b??????1?????1???11?1) z |= 4'b0010; 
	if(x==?20'b?????1??????1???11?1) z |= 4'b0010; 
	if(x==?20'b??????1????????111?1) z |= 4'b0001; 
	if(x==?20'b?????1?????????111?1) z |= 4'b0001; 
	if(x==?20'b1?????1?????????111?) z |= 4'b1000; 
	if(x==?20'b1????1??????????111?) z |= 4'b1000; 
	if(x==?20'b???1??1?????????111?) z |= 4'b0100; 
	if(x==?20'b???1?1??????????111?) z |= 4'b0100; 
	if(x==?20'b??????????1?1???111?) z |= 4'b0010; 
	if(x==?20'b?????????1??1???111?) z |= 4'b0010; 
	if(x==?20'b??????????1????1111?) z |= 4'b0001; 
	if(x==?20'b?????????1?????1111?) z |= 4'b0001; 
	if(x==?20'b?????1??1?1??????11?) z |= 4'b1010; 
	if(x==?20'b????1?1??1???????11?) z |= 4'b1010; 
	if(x==?20'b??????1??1?1?????11?) z |= 4'b0101; 
	if(x==?20'b?????1?1??1??????11?) z |= 4'b0101; 
	if(x==?20'b1???????????????1111) z |= 4'b1000; 
	if(x==?20'b???1????????????1111) z |= 4'b0100; 
	if(x==?20'b????????????1???1111) z |= 4'b0010; 
	if(x==?20'b???????????????11111) z |= 4'b0001; 
	if(x==?20'b??1???1???1?????11??) z |= 4'b1000; 
	if(x==?20'b?1???1???1??????11??) z |= 4'b0100; 
	if(x==?20'b??????1???1???1?11??) z |= 4'b0010; 
	if(x==?20'b?????1???1???1??11??) z |= 4'b0001; 
	if(x==?20'b?????11??11?????1?1?) z |= 4'b1111; 
	if(x==?20'b??1???????1?????11?1) z |= 4'b1000; 
	if(x==?20'b?1???????1??????11?1) z |= 4'b0100; 
	if(x==?20'b??????1???????1?11?1) z |= 4'b0010; 
	if(x==?20'b?????1???????1??11?1) z |= 4'b0001; 
	if(x==?20'b??1???1?????????111?) z |= 4'b1000; 
	if(x==?20'b?1???1??????????111?) z |= 4'b0100; 
	if(x==?20'b??????????1???1?111?) z |= 4'b0010; 
	if(x==?20'b?????????1???1??111?) z |= 4'b0001; 
	if(x==?20'b????????1???????1111) z |= 4'b1000; 
	if(x==?20'b???????????1????1111) z |= 4'b0100; 
	if(x==?20'b????1???????????1111) z |= 4'b0010; 
	if(x==?20'b???????1????????1111) z |= 4'b0001; 
	if(x==?20'b??1?????????????1111) z |= 4'b1000; 
	if(x==?20'b?1??????????????1111) z |= 4'b0100; 
	if(x==?20'b??????????????1?1111) z |= 4'b0010; 
	if(x==?20'b?????????????1??1111) z |= 4'b0001; 
	if(x==?20'b?????????11?????1?11) z |= 4'b1100; 
	if(x==?20'b?????11?????????1?11) z |= 4'b0011; 
	if(x==?20'b????1???1???????111?) z |= 4'b1010; 
	if(x==?20'b???????1???1????111?) z |= 4'b0101; 
	if(x==?20'b??????????1?????1111) z |= 4'b1000; 
	if(x==?20'b?????????1??????1111) z |= 4'b0100; 
	if(x==?20'b??????1?????????1111) z |= 4'b0010; 
	if(x==?20'b?????1??????????1111) z |= 4'b0001; 
	if(x==?20'b?1????1???1?????11??) z |= 4'b1100; 
	if(x==?20'b??1??1????1?????11??) z |= 4'b1100; 
	if(x==?20'b?1???1????1?????11??) z |= 4'b1100; 
	if(x==?20'b??1???1??1??????11??) z |= 4'b1100; 
	if(x==?20'b?1????1??1??????11??) z |= 4'b1100; 
	if(x==?20'b??1??1???1??????11??) z |= 4'b1100; 
	if(x==?20'b?????1????1???1?11??) z |= 4'b0011; 
	if(x==?20'b??????1??1????1?11??) z |= 4'b0011; 
	if(x==?20'b?????1???1????1?11??) z |= 4'b0011; 
	if(x==?20'b??????1???1??1??11??) z |= 4'b0011; 
	if(x==?20'b?????1????1??1??11??) z |= 4'b0011; 
	if(x==?20'b??????1??1???1??11??) z |= 4'b0011; 
	if(x==?20'b????11??????????1??1) z |= 4'b1000; 
	if(x==?20'b??????11????????1??1) z |= 4'b0100; 
	if(x==?20'b????????11??????1??1) z |= 4'b0010; 
	if(x==?20'b??????????11????1??1) z |= 4'b0001; 
	if(x==?20'b?1???1???1???????1??) z |= 4'b1000; 
	if(x==?20'b??1???1???1??????1??) z |= 4'b0100; 
	if(x==?20'b?????1???1???1???1??) z |= 4'b0010; 
	if(x==?20'b??????1???1???1??1??) z |= 4'b0001; 
	if(x==?20'b?1????????1?????11?1) z |= 4'b1100; 
	if(x==?20'b??1??????1??????11?1) z |= 4'b1100; 
	if(x==?20'b?????1????????1?11?1) z |= 4'b0011; 
	if(x==?20'b??????1??????1??11?1) z |= 4'b0011; 
	if(x==?20'b????1?????1?????111?) z |= 4'b1010; 
	if(x==?20'b????1????1??????111?) z |= 4'b1010; 
	if(x==?20'b??????1?1???????111?) z |= 4'b1010; 
	if(x==?20'b?????1??1???????111?) z |= 4'b1010; 
	if(x==?20'b??????1????1????111?) z |= 4'b0101; 
	if(x==?20'b?????1?????1????111?) z |= 4'b0101; 
	if(x==?20'b???????1??1?????111?) z |= 4'b0101; 
	if(x==?20'b???????1?1??????111?) z |= 4'b0101; 
	if(x==?20'b????1?1??????????1?1) z |= 4'b1000; 
	if(x==?20'b?????1?1?????????1?1) z |= 4'b0100; 
	if(x==?20'b????????1?1??????1?1) z |= 4'b0010; 
	if(x==?20'b?????????1?1?????1?1) z |= 4'b0001; 
	if(x==?20'b?1????1?????????111?) z |= 4'b1100; 
	if(x==?20'b??1??1??????????111?) z |= 4'b1100; 
	if(x==?20'b?????????1????1?111?) z |= 4'b0011; 
	if(x==?20'b??????????1??1??111?) z |= 4'b0011; 
	if(x==?20'b?1???????1???????1?1) z |= 4'b1000; 
	if(x==?20'b??1???????1??????1?1) z |= 4'b0100; 
	if(x==?20'b?????1???????1???1?1) z |= 4'b0010; 
	if(x==?20'b??????1???????1??1?1) z |= 4'b0001; 
	if(x==?20'b?1???1???????????11?) z |= 4'b1000; 
	if(x==?20'b??1???1??????????11?) z |= 4'b0100; 
	if(x==?20'b?????????1???1???11?) z |= 4'b0010; 
	if(x==?20'b??????????1???1??11?) z |= 4'b0001; 
	if(x==?20'b?1???????????????111) z |= 4'b1000; 
	if(x==?20'b??1??????????????111) z |= 4'b0100; 
	if(x==?20'b?????????????1???111) z |= 4'b0010; 
	if(x==?20'b??????????????1??111) z |= 4'b0001; 
	if(x==?20'b??????1???1?????111?) z |= 4'b1010; 
	if(x==?20'b?????1???1??????111?) z |= 4'b0101; 
	if(x==?20'b?????????1???????111) z |= 4'b1000; 
	if(x==?20'b??????????1??????111) z |= 4'b0100; 
	if(x==?20'b?????1???????????111) z |= 4'b0010; 
	if(x==?20'b??????1??????????111) z |= 4'b0001; 
	if(x==?20'b????1???????????11?1) z |= 4'b1000; 
	if(x==?20'b???????1????????11?1) z |= 4'b0100; 
	if(x==?20'b????????1???????11?1) z |= 4'b0010; 
	if(x==?20'b???????????1????11?1) z |= 4'b0001; 
	if(x==?20'b?????11?????????1??1) z |= 4'b1100; 
	if(x==?20'b?????????11?????1??1) z |= 4'b0011; 
	if(x==?20'b?????1???1???????11?) z |= 4'b1010; 
	if(x==?20'b??????1???1??????11?) z |= 4'b0101; 
	if(x==?20'b??????1?????????11?1) z |= 4'b1000; 
	if(x==?20'b?????1??????????11?1) z |= 4'b0100; 
	if(x==?20'b??????????1?????11?1) z |= 4'b0010; 
	if(x==?20'b?????????1??????11?1) z |= 4'b0001; 
	if(x==?20'b?????1????1?????111?) z |= 4'b1111; 
	if(x==?20'b??????1??1??????111?) z |= 4'b1111; 
	if(x==?20'b?????1???????????1?1) z |= 4'b1000; 
	if(x==?20'b??????1??????????1?1) z |= 4'b0100; 
	if(x==?20'b?????????1???????1?1) z |= 4'b0010; 
	if(x==?20'b??????????1??????1?1) z |= 4'b0001; 
end 
`endif
endmodule