module gb4_opt(
    input [19:0] x,
    output logic [3:0] z
);
always_comb begin 
	 z = 4'b0000;
	if(x==?20'b111?1???11??????000?) z |= 4'b1000; 
	if(x==?20'b111?1?1?1???????000?) z |= 4'b1000; 
	if(x==?20'b?111???1??11????000?) z |= 4'b0100; 
	if(x==?20'b?111?1?1???1????000?) z |= 4'b0100; 
	if(x==?20'b????1???1?1?111?000?) z |= 4'b0010; 
	if(x==?20'b????11??1???111?000?) z |= 4'b0010; 
	if(x==?20'b???????1?1?1?111000?) z |= 4'b0001; 
	if(x==?20'b??????11???1?111000?) z |= 4'b0001; 
	if(x==?20'b111?1???111??????00?) z |= 4'b1000; 
	if(x==?20'b111?1?1?1?1??????00?) z |= 4'b1000; 
	if(x==?20'b111?1?1?11??????0?0?) z |= 4'b1000; 
	if(x==?20'b?111???1?111?????00?) z |= 4'b0100; 
	if(x==?20'b?111?1?1?1?1?????00?) z |= 4'b0100; 
	if(x==?20'b?111?1?1??11????0?0?) z |= 4'b0100; 
	if(x==?20'b????1?1?1?1?111??00?) z |= 4'b0010; 
	if(x==?20'b????111?1???111??00?) z |= 4'b0010; 
	if(x==?20'b????11??1?1?111?0?0?) z |= 4'b0010; 
	if(x==?20'b?????1?1?1?1?111?00?) z |= 4'b0001; 
	if(x==?20'b?????111???1?111?00?) z |= 4'b0001; 
	if(x==?20'b??????11?1?1?1110?0?) z |= 4'b0001; 
	if(x==?20'b111?1?1?111???????0?) z |= 4'b1000; 
	if(x==?20'b111?11??11??????00??) z |= 4'b1000; 
	if(x==?20'b111?111?1???????00??) z |= 4'b1000; 
	if(x==?20'b?111?1?1?111??????0?) z |= 4'b0100; 
	if(x==?20'b?111??11??11????00??) z |= 4'b0100; 
	if(x==?20'b?111?111???1????00??) z |= 4'b0100; 
	if(x==?20'b????111?1?1?111???0?) z |= 4'b0010; 
	if(x==?20'b????1???111?111?00??) z |= 4'b0010; 
	if(x==?20'b????11??11??111?00??) z |= 4'b0010; 
	if(x==?20'b?????111?1?1?111??0?) z |= 4'b0001; 
	if(x==?20'b???????1?111?11100??) z |= 4'b0001; 
	if(x==?20'b??????11??11?11100??) z |= 4'b0001; 
	if(x==?20'b111?11??111??????0??) z |= 4'b1000; 
	if(x==?20'b111?111?1?1??????0??) z |= 4'b1000; 
	if(x==?20'b111?111?11??????0???) z |= 4'b1000; 
	if(x==?20'b?111??11?111?????0??) z |= 4'b0100; 
	if(x==?20'b?111?111?1?1?????0??) z |= 4'b0100; 
	if(x==?20'b?111?111??11????0???) z |= 4'b0100; 
	if(x==?20'b????1?1?111?111??0??) z |= 4'b0010; 
	if(x==?20'b????111?11??111??0??) z |= 4'b0010; 
	if(x==?20'b????11??111?111?0???) z |= 4'b0010; 
	if(x==?20'b?????1?1?111?111?0??) z |= 4'b0001; 
	if(x==?20'b?????111??11?111?0??) z |= 4'b0001; 
	if(x==?20'b??????11?111?1110???) z |= 4'b0001; 
	if(x==?20'b111?111?111?????????) z |= 4'b1000; 
	if(x==?20'b?111?111?111????????) z |= 4'b0100; 
	if(x==?20'b????111?111?111?????) z |= 4'b0010; 
	if(x==?20'b?????111?111?111????) z |= 4'b0001; 
	if(x==?20'b11??1???111?????000?) z |= 4'b1000; 
	if(x==?20'b111?1????11?????000?) z |= 4'b1000; 
	if(x==?20'b11??1?1?1?1?????000?) z |= 4'b1000; 
	if(x==?20'b111?1?1???1?????000?) z |= 4'b1000; 
	if(x==?20'b1?1?1?1?11??????000?) z |= 4'b1000; 
	if(x==?20'b111???1?11??????000?) z |= 4'b1000; 
	if(x==?20'b??11???1?111????000?) z |= 4'b0100; 
	if(x==?20'b?1?1?1?1??11????000?) z |= 4'b0100; 
	if(x==?20'b?111?1????11????000?) z |= 4'b0100; 
	if(x==?20'b??11?1?1?1?1????000?) z |= 4'b0100; 
	if(x==?20'b?111???1?11?????000?) z |= 4'b0100; 
	if(x==?20'b?111?1?1?1??????000?) z |= 4'b0100; 
	if(x==?20'b??????1?1?1?111?000?) z |= 4'b0010; 
	if(x==?20'b????11????1?111?000?) z |= 4'b0010; 
	if(x==?20'b?????11?1???111?000?) z |= 4'b0010; 
	if(x==?20'b????11??1?1?1?1?000?) z |= 4'b0010; 
	if(x==?20'b????1?1?1?1?11??000?) z |= 4'b0010; 
	if(x==?20'b????111?1???11??000?) z |= 4'b0010; 
	if(x==?20'b?????1???1?1?111000?) z |= 4'b0001; 
	if(x==?20'b?????11????1?111000?) z |= 4'b0001; 
	if(x==?20'b??????11?1???111000?) z |= 4'b0001; 
	if(x==?20'b?????1?1?1?1??11000?) z |= 4'b0001; 
	if(x==?20'b?????111???1??11000?) z |= 4'b0001; 
	if(x==?20'b??????11?1?1?1?1000?) z |= 4'b0001; 
	if(x==?20'b1?1?1?1?111??????00?) z |= 4'b1000; 
	if(x==?20'b111???1?111??????00?) z |= 4'b1000; 
	if(x==?20'b11??1?1?111?????0?0?) z |= 4'b1000; 
	if(x==?20'b111?1?1??11?????0?0?) z |= 4'b1000; 
	if(x==?20'b?1?1?1?1?111?????00?) z |= 4'b0100; 
	if(x==?20'b?111?1???111?????00?) z |= 4'b0100; 
	if(x==?20'b??11?1?1?111????0?0?) z |= 4'b0100; 
	if(x==?20'b?111?1?1?11?????0?0?) z |= 4'b0100; 
	if(x==?20'b????111???1?111??00?) z |= 4'b0010; 
	if(x==?20'b????111?1?1?1?1??00?) z |= 4'b0010; 
	if(x==?20'b?????11?1?1?111?0?0?) z |= 4'b0010; 
	if(x==?20'b????111?1?1?11??0?0?) z |= 4'b0010; 
	if(x==?20'b?????111?1???111?00?) z |= 4'b0001; 
	if(x==?20'b?????111?1?1?1?1?00?) z |= 4'b0001; 
	if(x==?20'b?????11??1?1?1110?0?) z |= 4'b0001; 
	if(x==?20'b?????111?1?1??110?0?) z |= 4'b0001; 
	if(x==?20'b11??11??111?????00??) z |= 4'b1000; 
	if(x==?20'b111?11???11?????00??) z |= 4'b1000; 
	if(x==?20'b11??111?1?1?????00??) z |= 4'b1000; 
	if(x==?20'b111?111???1?????00??) z |= 4'b1000; 
	if(x==?20'b1?1?111?11??????00??) z |= 4'b1000; 
	if(x==?20'b111??11?11??????00??) z |= 4'b1000; 
	if(x==?20'b??11??11?111????00??) z |= 4'b0100; 
	if(x==?20'b?1?1?111??11????00??) z |= 4'b0100; 
	if(x==?20'b?111?11???11????00??) z |= 4'b0100; 
	if(x==?20'b??11?111?1?1????00??) z |= 4'b0100; 
	if(x==?20'b?111??11?11?????00??) z |= 4'b0100; 
	if(x==?20'b?111?111?1??????00??) z |= 4'b0100; 
	if(x==?20'b??????1?111?111?00??) z |= 4'b0010; 
	if(x==?20'b????11???11?111?00??) z |= 4'b0010; 
	if(x==?20'b?????11?11??111?00??) z |= 4'b0010; 
	if(x==?20'b????11??111?1?1?00??) z |= 4'b0010; 
	if(x==?20'b????1?1?111?11??00??) z |= 4'b0010; 
	if(x==?20'b????111?11??11??00??) z |= 4'b0010; 
	if(x==?20'b?????1???111?11100??) z |= 4'b0001; 
	if(x==?20'b?????11???11?11100??) z |= 4'b0001; 
	if(x==?20'b??????11?11??11100??) z |= 4'b0001; 
	if(x==?20'b?????1?1?111??1100??) z |= 4'b0001; 
	if(x==?20'b?????111??11??1100??) z |= 4'b0001; 
	if(x==?20'b??????11?111?1?100??) z |= 4'b0001; 
	if(x==?20'b1?1?111?111??????0??) z |= 4'b1000; 
	if(x==?20'b111??11?111??????0??) z |= 4'b1000; 
	if(x==?20'b11??111?111?????0???) z |= 4'b1000; 
	if(x==?20'b111?111??11?????0???) z |= 4'b1000; 
	if(x==?20'b?1?1?111?111?????0??) z |= 4'b0100; 
	if(x==?20'b?111?11??111?????0??) z |= 4'b0100; 
	if(x==?20'b??11?111?111????0???) z |= 4'b0100; 
	if(x==?20'b?111?111?11?????0???) z |= 4'b0100; 
	if(x==?20'b????111??11?111??0??) z |= 4'b0010; 
	if(x==?20'b????111?111?1?1??0??) z |= 4'b0010; 
	if(x==?20'b?????11?111?111?0???) z |= 4'b0010; 
	if(x==?20'b????111?111?11??0???) z |= 4'b0010; 
	if(x==?20'b?????111?11??111?0??) z |= 4'b0001; 
	if(x==?20'b?????111?111?1?1?0??) z |= 4'b0001; 
	if(x==?20'b?????11??111?1110???) z |= 4'b0001; 
	if(x==?20'b?????111?111??110???) z |= 4'b0001; 
	if(x==?20'b?11?1???111?????000?) z |= 4'b1000; 
	if(x==?20'b?11?1?1?1?1?????000?) z |= 4'b1000; 
	if(x==?20'b?11????1?111????000?) z |= 4'b0100; 
	if(x==?20'b?11??1?1?1?1????000?) z |= 4'b0100; 
	if(x==?20'b????1?1?1?1??11?000?) z |= 4'b0010; 
	if(x==?20'b????111?1????11?000?) z |= 4'b0010; 
	if(x==?20'b?????1?1?1?1?11?000?) z |= 4'b0001; 
	if(x==?20'b?????111???1?11?000?) z |= 4'b0001; 
	if(x==?20'b?11?1?1?111?????0?0?) z |= 4'b1000; 
	if(x==?20'b?11??1?1?111????0?0?) z |= 4'b0100; 
	if(x==?20'b????111?1?1??11?0?0?) z |= 4'b0010; 
	if(x==?20'b?????111?1?1?11?0?0?) z |= 4'b0001; 
	if(x==?20'b?11?11??111?????00??) z |= 4'b1000; 
	if(x==?20'b?11?111?1?1?????00??) z |= 4'b1000; 
	if(x==?20'b?11???11?111????00??) z |= 4'b0100; 
	if(x==?20'b?11??111?1?1????00??) z |= 4'b0100; 
	if(x==?20'b????1?1?111??11?00??) z |= 4'b0010; 
	if(x==?20'b????111?11???11?00??) z |= 4'b0010; 
	if(x==?20'b?????1?1?111?11?00??) z |= 4'b0001; 
	if(x==?20'b?????111??11?11?00??) z |= 4'b0001; 
	if(x==?20'b?11?111?111?????0???) z |= 4'b1000; 
	if(x==?20'b?11??111?111????0???) z |= 4'b0100; 
	if(x==?20'b????111?111??11?0???) z |= 4'b0010; 
	if(x==?20'b?????111?111?11?0???) z |= 4'b0001; 
	if(x==?20'b1???1?1?111?????000?) z |= 4'b1000; 
	if(x==?20'b11????1?111?????000?) z |= 4'b1000; 
	if(x==?20'b1?1?1?1??11?????000?) z |= 4'b1000; 
	if(x==?20'b111???1??11?????000?) z |= 4'b1000; 
	if(x==?20'b???1?1?1?111????000?) z |= 4'b0100; 
	if(x==?20'b??11?1???111????000?) z |= 4'b0100; 
	if(x==?20'b?1?1?1?1?11?????000?) z |= 4'b0100; 
	if(x==?20'b?111?1???11?????000?) z |= 4'b0100; 
	if(x==?20'b?????11???1?111?000?) z |= 4'b0010; 
	if(x==?20'b?????11?1?1?1?1?000?) z |= 4'b0010; 
	if(x==?20'b????111???1?11??000?) z |= 4'b0010; 
	if(x==?20'b????111?1?1?1???000?) z |= 4'b0010; 
	if(x==?20'b?????11??1???111000?) z |= 4'b0001; 
	if(x==?20'b?????111?1????11000?) z |= 4'b0001; 
	if(x==?20'b?????11??1?1?1?1000?) z |= 4'b0001; 
	if(x==?20'b?????111?1?1???1000?) z |= 4'b0001; 
	if(x==?20'b1???111?111?????00??) z |= 4'b1000; 
	if(x==?20'b11???11?111?????00??) z |= 4'b1000; 
	if(x==?20'b1?1?111??11?????00??) z |= 4'b1000; 
	if(x==?20'b111??11??11?????00??) z |= 4'b1000; 
	if(x==?20'b???1?111?111????00??) z |= 4'b0100; 
	if(x==?20'b??11?11??111????00??) z |= 4'b0100; 
	if(x==?20'b?1?1?111?11?????00??) z |= 4'b0100; 
	if(x==?20'b?111?11??11?????00??) z |= 4'b0100; 
	if(x==?20'b?????11??11?111?00??) z |= 4'b0010; 
	if(x==?20'b?????11?111?1?1?00??) z |= 4'b0010; 
	if(x==?20'b????111??11?11??00??) z |= 4'b0010; 
	if(x==?20'b????111?111?1???00??) z |= 4'b0010; 
	if(x==?20'b?????11??11??11100??) z |= 4'b0001; 
	if(x==?20'b?????111?11???1100??) z |= 4'b0001; 
	if(x==?20'b?????11??111?1?100??) z |= 4'b0001; 
	if(x==?20'b?????111?111???100??) z |= 4'b0001; 
	if(x==?20'b111?11??1???????0?0?) z |= 4'b1000; 
	if(x==?20'b?111??11???1????0?0?) z |= 4'b0100; 
	if(x==?20'b????1???11??111?0?0?) z |= 4'b0010; 
	if(x==?20'b???????1??11?1110?0?) z |= 4'b0001; 
	if(x==?20'b111?11??1?1???????0?) z |= 4'b1000; 
	if(x==?20'b?111??11?1?1??????0?) z |= 4'b0100; 
	if(x==?20'b????1?1?11??111???0?) z |= 4'b0010; 
	if(x==?20'b?????1?1??11?111??0?) z |= 4'b0001; 
	if(x==?20'b??1?1?1?111?????000?) z |= 4'b1000; 
	if(x==?20'b?11???1?111?????000?) z |= 4'b1000; 
	if(x==?20'b?1???1?1?111????000?) z |= 4'b0100; 
	if(x==?20'b?11??1???111????000?) z |= 4'b0100; 
	if(x==?20'b????111???1??11?000?) z |= 4'b0010; 
	if(x==?20'b????111?1?1???1?000?) z |= 4'b0010; 
	if(x==?20'b?????111?1???11?000?) z |= 4'b0001; 
	if(x==?20'b?????111?1?1?1??000?) z |= 4'b0001; 
	if(x==?20'b??1?111?111?????00??) z |= 4'b1000; 
	if(x==?20'b?11??11?111?????00??) z |= 4'b1000; 
	if(x==?20'b?1???111?111????00??) z |= 4'b0100; 
	if(x==?20'b?11??11??111????00??) z |= 4'b0100; 
	if(x==?20'b????111??11??11?00??) z |= 4'b0010; 
	if(x==?20'b????111?111???1?00??) z |= 4'b0010; 
	if(x==?20'b?????111?11??11?00??) z |= 4'b0001; 
	if(x==?20'b?????111?111?1??00??) z |= 4'b0001; 
	if(x==?20'b1?1?11??1???????000?) z |= 4'b1000; 
	if(x==?20'b111??1??1???????000?) z |= 4'b1000; 
	if(x==?20'b?1?1??11???1????000?) z |= 4'b0100; 
	if(x==?20'b?111??1????1????000?) z |= 4'b0100; 
	if(x==?20'b????1????1??111?000?) z |= 4'b0010; 
	if(x==?20'b????1???11??1?1?000?) z |= 4'b0010; 
	if(x==?20'b???????1??1??111000?) z |= 4'b0001; 
	if(x==?20'b???????1??11?1?1000?) z |= 4'b0001; 
	if(x==?20'b1?1?11??1?1??????00?) z |= 4'b1000; 
	if(x==?20'b111??1??1?1??????00?) z |= 4'b1000; 
	if(x==?20'b11??1?1?11???????00?) z |= 4'b1000; 
	if(x==?20'b111?1?1??1???????00?) z |= 4'b1000; 
	if(x==?20'b11??11??1?1?????0?0?) z |= 4'b1000; 
	if(x==?20'b111?11????1?????0?0?) z |= 4'b1000; 
	if(x==?20'b1?1?11??11??????0?0?) z |= 4'b1000; 
	if(x==?20'b111??1??11??????0?0?) z |= 4'b1000; 
	if(x==?20'b1?1?111?1???????0?0?) z |= 4'b1000; 
	if(x==?20'b111??11?1???????0?0?) z |= 4'b1000; 
	if(x==?20'b??11?1?1??11?????00?) z |= 4'b0100; 
	if(x==?20'b?1?1??11?1?1?????00?) z |= 4'b0100; 
	if(x==?20'b?111??1??1?1?????00?) z |= 4'b0100; 
	if(x==?20'b?111?1?1??1??????00?) z |= 4'b0100; 
	if(x==?20'b?1?1??11??11????0?0?) z |= 4'b0100; 
	if(x==?20'b?111??1???11????0?0?) z |= 4'b0100; 
	if(x==?20'b??11??11?1?1????0?0?) z |= 4'b0100; 
	if(x==?20'b?1?1?111???1????0?0?) z |= 4'b0100; 
	if(x==?20'b?111?11????1????0?0?) z |= 4'b0100; 
	if(x==?20'b?111??11?1??????0?0?) z |= 4'b0100; 
	if(x==?20'b?????1??1?1?111??00?) z |= 4'b0010; 
	if(x==?20'b????1?1??1??111??00?) z |= 4'b0010; 
	if(x==?20'b????1?1?11??1?1??00?) z |= 4'b0010; 
	if(x==?20'b????11??1?1?11???00?) z |= 4'b0010; 
	if(x==?20'b????1????11?111?0?0?) z |= 4'b0010; 
	if(x==?20'b??????1?11??111?0?0?) z |= 4'b0010; 
	if(x==?20'b????11???1??111?0?0?) z |= 4'b0010; 
	if(x==?20'b????1???111?1?1?0?0?) z |= 4'b0010; 
	if(x==?20'b????11??11??1?1?0?0?) z |= 4'b0010; 
	if(x==?20'b????1?1?11??11??0?0?) z |= 4'b0010; 
	if(x==?20'b??????1??1?1?111?00?) z |= 4'b0001; 
	if(x==?20'b?????1?1??1??111?00?) z |= 4'b0001; 
	if(x==?20'b??????11?1?1??11?00?) z |= 4'b0001; 
	if(x==?20'b?????1?1??11?1?1?00?) z |= 4'b0001; 
	if(x==?20'b?????1????11?1110?0?) z |= 4'b0001; 
	if(x==?20'b???????1?11??1110?0?) z |= 4'b0001; 
	if(x==?20'b??????11??1??1110?0?) z |= 4'b0001; 
	if(x==?20'b?????1?1??11??110?0?) z |= 4'b0001; 
	if(x==?20'b???????1?111?1?10?0?) z |= 4'b0001; 
	if(x==?20'b??????11??11?1?10?0?) z |= 4'b0001; 
	if(x==?20'b1?1?11??111???????0?) z |= 4'b1000; 
	if(x==?20'b111??1??111???????0?) z |= 4'b1000; 
	if(x==?20'b1?1?111?1?1???????0?) z |= 4'b1000; 
	if(x==?20'b111??11?1?1???????0?) z |= 4'b1000; 
	if(x==?20'b?1?1??11?111??????0?) z |= 4'b0100; 
	if(x==?20'b?111??1??111??????0?) z |= 4'b0100; 
	if(x==?20'b?1?1?111?1?1??????0?) z |= 4'b0100; 
	if(x==?20'b?111?11??1?1??????0?) z |= 4'b0100; 
	if(x==?20'b????1?1??11?111???0?) z |= 4'b0010; 
	if(x==?20'b????111??1??111???0?) z |= 4'b0010; 
	if(x==?20'b????1?1?111?1?1???0?) z |= 4'b0010; 
	if(x==?20'b????111?11??1?1???0?) z |= 4'b0010; 
	if(x==?20'b?????1?1?11??111??0?) z |= 4'b0001; 
	if(x==?20'b?????111??1??111??0?) z |= 4'b0001; 
	if(x==?20'b?????1?1?111?1?1??0?) z |= 4'b0001; 
	if(x==?20'b?????111??11?1?1??0?) z |= 4'b0001; 
	if(x==?20'b11??111?11???????0??) z |= 4'b1000; 
	if(x==?20'b111?111??1???????0??) z |= 4'b1000; 
	if(x==?20'b??11?111??11?????0??) z |= 4'b0100; 
	if(x==?20'b?111?111??1??????0??) z |= 4'b0100; 
	if(x==?20'b?????1??111?111??0??) z |= 4'b0010; 
	if(x==?20'b????11??111?11???0??) z |= 4'b0010; 
	if(x==?20'b??????1??111?111?0??) z |= 4'b0001; 
	if(x==?20'b??????11?111??11?0??) z |= 4'b0001; 
	if(x==?20'b?11?1?1?11???????00?) z |= 4'b1000; 
	if(x==?20'b?11?11??1?1?????0?0?) z |= 4'b1000; 
	if(x==?20'b?11??1?1??11?????00?) z |= 4'b0100; 
	if(x==?20'b?11???11?1?1????0?0?) z |= 4'b0100; 
	if(x==?20'b????11??1?1??11??00?) z |= 4'b0010; 
	if(x==?20'b????1?1?11???11?0?0?) z |= 4'b0010; 
	if(x==?20'b??????11?1?1?11??00?) z |= 4'b0001; 
	if(x==?20'b?????1?1??11?11?0?0?) z |= 4'b0001; 
	if(x==?20'b?11?111?11???????0??) z |= 4'b1000; 
	if(x==?20'b?11??111??11?????0??) z |= 4'b0100; 
	if(x==?20'b????11??111??11??0??) z |= 4'b0010; 
	if(x==?20'b??????11?111?11??0??) z |= 4'b0001; 
	if(x==?20'b1???11??1?1?????000?) z |= 4'b1000; 
	if(x==?20'b11???1??1?1?????000?) z |= 4'b1000; 
	if(x==?20'b1?1?11????1?????000?) z |= 4'b1000; 
	if(x==?20'b111??1????1?????000?) z |= 4'b1000; 
	if(x==?20'b1?1??1??11??????000?) z |= 4'b1000; 
	if(x==?20'b11??1?1??1??????000?) z |= 4'b1000; 
	if(x==?20'b1?1??11?1???????000?) z |= 4'b1000; 
	if(x==?20'b?1?1??1???11????000?) z |= 4'b0100; 
	if(x==?20'b???1??11?1?1????000?) z |= 4'b0100; 
	if(x==?20'b??11??1??1?1????000?) z |= 4'b0100; 
	if(x==?20'b?1?1?11????1????000?) z |= 4'b0100; 
	if(x==?20'b??11?1?1??1?????000?) z |= 4'b0100; 
	if(x==?20'b?1?1??11?1??????000?) z |= 4'b0100; 
	if(x==?20'b?111??1??1??????000?) z |= 4'b0100; 
	if(x==?20'b??????1??1??111?000?) z |= 4'b0010; 
	if(x==?20'b????1????11?1?1?000?) z |= 4'b0010; 
	if(x==?20'b??????1?11??1?1?000?) z |= 4'b0010; 
	if(x==?20'b????11???1??1?1?000?) z |= 4'b0010; 
	if(x==?20'b?????1??1?1?11??000?) z |= 4'b0010; 
	if(x==?20'b????1?1??1??11??000?) z |= 4'b0010; 
	if(x==?20'b????1?1?11??1???000?) z |= 4'b0010; 
	if(x==?20'b?????1????1??111000?) z |= 4'b0001; 
	if(x==?20'b??????1??1?1??11000?) z |= 4'b0001; 
	if(x==?20'b?????1?1??1???11000?) z |= 4'b0001; 
	if(x==?20'b?????1????11?1?1000?) z |= 4'b0001; 
	if(x==?20'b???????1?11??1?1000?) z |= 4'b0001; 
	if(x==?20'b??????11??1??1?1000?) z |= 4'b0001; 
	if(x==?20'b?????1?1??11???1000?) z |= 4'b0001; 
	if(x==?20'b1?1??1??111??????00?) z |= 4'b1000; 
	if(x==?20'b11??1?1??11??????00?) z |= 4'b1000; 
	if(x==?20'b1?1??11?1?1??????00?) z |= 4'b1000; 
	if(x==?20'b1???11??111?????0?0?) z |= 4'b1000; 
	if(x==?20'b11???1??111?????0?0?) z |= 4'b1000; 
	if(x==?20'b1?1?11???11?????0?0?) z |= 4'b1000; 
	if(x==?20'b111??1???11?????0?0?) z |= 4'b1000; 
	if(x==?20'b1???111?1?1?????0?0?) z |= 4'b1000; 
	if(x==?20'b11???11?1?1?????0?0?) z |= 4'b1000; 
	if(x==?20'b1?1?111???1?????0?0?) z |= 4'b1000; 
	if(x==?20'b111??11???1?????0?0?) z |= 4'b1000; 
	if(x==?20'b1?1??11?11??????0?0?) z |= 4'b1000; 
	if(x==?20'b?1?1??1??111?????00?) z |= 4'b0100; 
	if(x==?20'b?1?1?11??1?1?????00?) z |= 4'b0100; 
	if(x==?20'b??11?1?1?11??????00?) z |= 4'b0100; 
	if(x==?20'b???1??11?111????0?0?) z |= 4'b0100; 
	if(x==?20'b??11??1??111????0?0?) z |= 4'b0100; 
	if(x==?20'b?1?1?11???11????0?0?) z |= 4'b0100; 
	if(x==?20'b???1?111?1?1????0?0?) z |= 4'b0100; 
	if(x==?20'b??11?11??1?1????0?0?) z |= 4'b0100; 
	if(x==?20'b?1?1??11?11?????0?0?) z |= 4'b0100; 
	if(x==?20'b?111??1??11?????0?0?) z |= 4'b0100; 
	if(x==?20'b?1?1?111?1??????0?0?) z |= 4'b0100; 
	if(x==?20'b?111?11??1??????0?0?) z |= 4'b0100; 
	if(x==?20'b????1?1??11?1?1??00?) z |= 4'b0010; 
	if(x==?20'b????111??1??1?1??00?) z |= 4'b0010; 
	if(x==?20'b?????11?1?1?11???00?) z |= 4'b0010; 
	if(x==?20'b??????1??11?111?0?0?) z |= 4'b0010; 
	if(x==?20'b?????11??1??111?0?0?) z |= 4'b0010; 
	if(x==?20'b??????1?111?1?1?0?0?) z |= 4'b0010; 
	if(x==?20'b????11???11?1?1?0?0?) z |= 4'b0010; 
	if(x==?20'b?????11?11??1?1?0?0?) z |= 4'b0010; 
	if(x==?20'b????1?1??11?11??0?0?) z |= 4'b0010; 
	if(x==?20'b????111??1??11??0?0?) z |= 4'b0010; 
	if(x==?20'b????1?1?111?1???0?0?) z |= 4'b0010; 
	if(x==?20'b????111?11??1???0?0?) z |= 4'b0010; 
	if(x==?20'b?????11??1?1??11?00?) z |= 4'b0001; 
	if(x==?20'b?????1?1?11??1?1?00?) z |= 4'b0001; 
	if(x==?20'b?????111??1??1?1?00?) z |= 4'b0001; 
	if(x==?20'b?????1???11??1110?0?) z |= 4'b0001; 
	if(x==?20'b?????11???1??1110?0?) z |= 4'b0001; 
	if(x==?20'b?????1?1?11???110?0?) z |= 4'b0001; 
	if(x==?20'b?????111??1???110?0?) z |= 4'b0001; 
	if(x==?20'b?????1???111?1?10?0?) z |= 4'b0001; 
	if(x==?20'b?????11???11?1?10?0?) z |= 4'b0001; 
	if(x==?20'b??????11?11??1?10?0?) z |= 4'b0001; 
	if(x==?20'b?????1?1?111???10?0?) z |= 4'b0001; 
	if(x==?20'b?????111??11???10?0?) z |= 4'b0001; 
	if(x==?20'b1?1??11?111???????0?) z |= 4'b1000; 
	if(x==?20'b11??111??1??????00??) z |= 4'b1000; 
	if(x==?20'b?1?1?11??111??????0?) z |= 4'b0100; 
	if(x==?20'b??11?111??1?????00??) z |= 4'b0100; 
	if(x==?20'b????111??11?1?1???0?) z |= 4'b0010; 
	if(x==?20'b?????1??111?11??00??) z |= 4'b0010; 
	if(x==?20'b?????111?11??1?1??0?) z |= 4'b0001; 
	if(x==?20'b??????1??111??1100??) z |= 4'b0001; 
	if(x==?20'b11??111??11??????0??) z |= 4'b1000; 
	if(x==?20'b??11?111?11??????0??) z |= 4'b0100; 
	if(x==?20'b?????11?111?11???0??) z |= 4'b0010; 
	if(x==?20'b?????11??111??11?0??) z |= 4'b0001; 
	if(x==?20'b111?1???1???????0??0) z |= 4'b1000; 
	if(x==?20'b?111???1???1????0??0) z |= 4'b0100; 
	if(x==?20'b????1???1???111?0??0) z |= 4'b0010; 
	if(x==?20'b???????1???1?1110??0) z |= 4'b0001; 
	if(x==?20'b111?1???1?1????????0) z |= 4'b1000; 
	if(x==?20'b?111???1?1?1???????0) z |= 4'b0100; 
	if(x==?20'b????1?1?1???111????0) z |= 4'b0010; 
	if(x==?20'b?????1?1???1?111???0) z |= 4'b0001; 
	if(x==?20'b??1?11??1?1?????000?) z |= 4'b1000; 
	if(x==?20'b?11??1??1?1?????000?) z |= 4'b1000; 
	if(x==?20'b?1??1?1?11??????000?) z |= 4'b1000; 
	if(x==?20'b?11?1?1??1??????000?) z |= 4'b1000; 
	if(x==?20'b??1??1?1??11????000?) z |= 4'b0100; 
	if(x==?20'b?1????11?1?1????000?) z |= 4'b0100; 
	if(x==?20'b?11???1??1?1????000?) z |= 4'b0100; 
	if(x==?20'b?11??1?1??1?????000?) z |= 4'b0100; 
	if(x==?20'b?????1??1?1??11?000?) z |= 4'b0010; 
	if(x==?20'b????1?1??1???11?000?) z |= 4'b0010; 
	if(x==?20'b????1?1?11????1?000?) z |= 4'b0010; 
	if(x==?20'b????11??1?1??1??000?) z |= 4'b0010; 
	if(x==?20'b??????1??1?1?11?000?) z |= 4'b0001; 
	if(x==?20'b?????1?1??1??11?000?) z |= 4'b0001; 
	if(x==?20'b??????11?1?1??1?000?) z |= 4'b0001; 
	if(x==?20'b?????1?1??11?1??000?) z |= 4'b0001; 
	if(x==?20'b?1??1?1?111??????00?) z |= 4'b1000; 
	if(x==?20'b?11?1?1??11??????00?) z |= 4'b1000; 
	if(x==?20'b??1?11??111?????0?0?) z |= 4'b1000; 
	if(x==?20'b?11??1??111?????0?0?) z |= 4'b1000; 
	if(x==?20'b??1?111?1?1?????0?0?) z |= 4'b1000; 
	if(x==?20'b?11??11?1?1?????0?0?) z |= 4'b1000; 
	if(x==?20'b??1??1?1?111?????00?) z |= 4'b0100; 
	if(x==?20'b?11??1?1?11??????00?) z |= 4'b0100; 
	if(x==?20'b?1????11?111????0?0?) z |= 4'b0100; 
	if(x==?20'b?11???1??111????0?0?) z |= 4'b0100; 
	if(x==?20'b?1???111?1?1????0?0?) z |= 4'b0100; 
	if(x==?20'b?11??11??1?1????0?0?) z |= 4'b0100; 
	if(x==?20'b?????11?1?1??11??00?) z |= 4'b0010; 
	if(x==?20'b????111?1?1??1???00?) z |= 4'b0010; 
	if(x==?20'b????1?1??11??11?0?0?) z |= 4'b0010; 
	if(x==?20'b????111??1???11?0?0?) z |= 4'b0010; 
	if(x==?20'b????1?1?111???1?0?0?) z |= 4'b0010; 
	if(x==?20'b????111?11????1?0?0?) z |= 4'b0010; 
	if(x==?20'b?????11??1?1?11??00?) z |= 4'b0001; 
	if(x==?20'b?????111?1?1??1??00?) z |= 4'b0001; 
	if(x==?20'b?????1?1?11??11?0?0?) z |= 4'b0001; 
	if(x==?20'b?????111??1??11?0?0?) z |= 4'b0001; 
	if(x==?20'b?????1?1?111?1??0?0?) z |= 4'b0001; 
	if(x==?20'b?????111??11?1??0?0?) z |= 4'b0001; 
	if(x==?20'b?1??111?11??????00??) z |= 4'b1000; 
	if(x==?20'b?11?111??1??????00??) z |= 4'b1000; 
	if(x==?20'b??1??111??11????00??) z |= 4'b0100; 
	if(x==?20'b?11??111??1?????00??) z |= 4'b0100; 
	if(x==?20'b?????1??111??11?00??) z |= 4'b0010; 
	if(x==?20'b????11??111??1??00??) z |= 4'b0010; 
	if(x==?20'b??????1??111?11?00??) z |= 4'b0001; 
	if(x==?20'b??????11?111??1?00??) z |= 4'b0001; 
	if(x==?20'b?1??111?111??????0??) z |= 4'b1000; 
	if(x==?20'b?11?111??11??????0??) z |= 4'b1000; 
	if(x==?20'b??1??111?111?????0??) z |= 4'b0100; 
	if(x==?20'b?11??111?11??????0??) z |= 4'b0100; 
	if(x==?20'b?????11?111??11??0??) z |= 4'b0010; 
	if(x==?20'b????111?111??1???0??) z |= 4'b0010; 
	if(x==?20'b?????11??111?11??0??) z |= 4'b0001; 
	if(x==?20'b?????111?111??1??0??) z |= 4'b0001; 
	if(x==?20'b1????1??111?????000?) z |= 4'b1000; 
	if(x==?20'b1?1??1???11?????000?) z |= 4'b1000; 
	if(x==?20'b1????11?1?1?????000?) z |= 4'b1000; 
	if(x==?20'b1?1??11???1?????000?) z |= 4'b1000; 
	if(x==?20'b???1??1??111????000?) z |= 4'b0100; 
	if(x==?20'b???1?11??1?1????000?) z |= 4'b0100; 
	if(x==?20'b?1?1??1??11?????000?) z |= 4'b0100; 
	if(x==?20'b?1?1?11??1??????000?) z |= 4'b0100; 
	if(x==?20'b??????1??11?1?1?000?) z |= 4'b0010; 
	if(x==?20'b?????11??1??1?1?000?) z |= 4'b0010; 
	if(x==?20'b????1?1??11?1???000?) z |= 4'b0010; 
	if(x==?20'b????111??1??1???000?) z |= 4'b0010; 
	if(x==?20'b?????1???11??1?1000?) z |= 4'b0001; 
	if(x==?20'b?????11???1??1?1000?) z |= 4'b0001; 
	if(x==?20'b?????1?1?11????1000?) z |= 4'b0001; 
	if(x==?20'b?????111??1????1000?) z |= 4'b0001; 
	if(x==?20'b1????11?111?????0?0?) z |= 4'b1000; 
	if(x==?20'b1?1??11??11?????0?0?) z |= 4'b1000; 
	if(x==?20'b???1?11??111????0?0?) z |= 4'b0100; 
	if(x==?20'b?1?1?11??11?????0?0?) z |= 4'b0100; 
	if(x==?20'b?????11??11?1?1?0?0?) z |= 4'b0010; 
	if(x==?20'b????111??11?1???0?0?) z |= 4'b0010; 
	if(x==?20'b?????11??11??1?10?0?) z |= 4'b0001; 
	if(x==?20'b?????111?11????10?0?) z |= 4'b0001; 
	if(x==?20'b11??11??1????????00?) z |= 4'b1000; 
	if(x==?20'b111?11???????????00?) z |= 4'b1000; 
	if(x==?20'b??11??11???1?????00?) z |= 4'b0100; 
	if(x==?20'b?111??11?????????00?) z |= 4'b0100; 
	if(x==?20'b????????11??111??00?) z |= 4'b0010; 
	if(x==?20'b????1???11??11???00?) z |= 4'b0010; 
	if(x==?20'b??????????11?111?00?) z |= 4'b0001; 
	if(x==?20'b???????1??11??11?00?) z |= 4'b0001; 
	if(x==?20'b11??11??11????????0?) z |= 4'b1000; 
	if(x==?20'b111?11???1????????0?) z |= 4'b1000; 
	if(x==?20'b11??111?1?????????0?) z |= 4'b1000; 
	if(x==?20'b111?111???????????0?) z |= 4'b1000; 
	if(x==?20'b??11??11??11??????0?) z |= 4'b0100; 
	if(x==?20'b??11?111???1??????0?) z |= 4'b0100; 
	if(x==?20'b?111??11??1???????0?) z |= 4'b0100; 
	if(x==?20'b?111?111??????????0?) z |= 4'b0100; 
	if(x==?20'b????????111?111???0?) z |= 4'b0010; 
	if(x==?20'b?????1??11??111???0?) z |= 4'b0010; 
	if(x==?20'b????1???111?11????0?) z |= 4'b0010; 
	if(x==?20'b????11??11??11????0?) z |= 4'b0010; 
	if(x==?20'b?????????111?111??0?) z |= 4'b0001; 
	if(x==?20'b??????1???11?111??0?) z |= 4'b0001; 
	if(x==?20'b???????1?111??11??0?) z |= 4'b0001; 
	if(x==?20'b??????11??11??11??0?) z |= 4'b0001; 
	if(x==?20'b1?1?1???1???????00?0) z |= 4'b1000; 
	if(x==?20'b111?????1???????00?0) z |= 4'b1000; 
	if(x==?20'b?1?1???1???1????00?0) z |= 4'b0100; 
	if(x==?20'b?111???????1????00?0) z |= 4'b0100; 
	if(x==?20'b????1???????111?00?0) z |= 4'b0010; 
	if(x==?20'b????1???1???1?1?00?0) z |= 4'b0010; 
	if(x==?20'b???????1?????11100?0) z |= 4'b0001; 
	if(x==?20'b???????1???1?1?100?0) z |= 4'b0001; 
	if(x==?20'b1?1?1???1?1??????0?0) z |= 4'b1000; 
	if(x==?20'b111?????1?1??????0?0) z |= 4'b1000; 
	if(x==?20'b11??1???1?1?????0??0) z |= 4'b1000; 
	if(x==?20'b111?1?????1?????0??0) z |= 4'b1000; 
	if(x==?20'b1?1?1???11??????0??0) z |= 4'b1000; 
	if(x==?20'b111?????11??????0??0) z |= 4'b1000; 
	if(x==?20'b1?1?1?1?1???????0??0) z |= 4'b1000; 
	if(x==?20'b111???1?1???????0??0) z |= 4'b1000; 
	if(x==?20'b?1?1???1?1?1?????0?0) z |= 4'b0100; 
	if(x==?20'b?111?????1?1?????0?0) z |= 4'b0100; 
	if(x==?20'b?1?1???1??11????0??0) z |= 4'b0100; 
	if(x==?20'b?111??????11????0??0) z |= 4'b0100; 
	if(x==?20'b??11???1?1?1????0??0) z |= 4'b0100; 
	if(x==?20'b?1?1?1?1???1????0??0) z |= 4'b0100; 
	if(x==?20'b?111?1?????1????0??0) z |= 4'b0100; 
	if(x==?20'b?111???1?1??????0??0) z |= 4'b0100; 
	if(x==?20'b????1?1?????111??0?0) z |= 4'b0010; 
	if(x==?20'b????1?1?1???1?1??0?0) z |= 4'b0010; 
	if(x==?20'b????1?????1?111?0??0) z |= 4'b0010; 
	if(x==?20'b??????1?1???111?0??0) z |= 4'b0010; 
	if(x==?20'b????11??????111?0??0) z |= 4'b0010; 
	if(x==?20'b????1???1?1?1?1?0??0) z |= 4'b0010; 
	if(x==?20'b????11??1???1?1?0??0) z |= 4'b0010; 
	if(x==?20'b????1?1?1???11??0??0) z |= 4'b0010; 
	if(x==?20'b?????1?1?????111?0?0) z |= 4'b0001; 
	if(x==?20'b?????1?1???1?1?1?0?0) z |= 4'b0001; 
	if(x==?20'b?????1?????1?1110??0) z |= 4'b0001; 
	if(x==?20'b???????1?1???1110??0) z |= 4'b0001; 
	if(x==?20'b??????11?????1110??0) z |= 4'b0001; 
	if(x==?20'b?????1?1???1??110??0) z |= 4'b0001; 
	if(x==?20'b???????1?1?1?1?10??0) z |= 4'b0001; 
	if(x==?20'b??????11???1?1?10??0) z |= 4'b0001; 
	if(x==?20'b1?1?1???111????????0) z |= 4'b1000; 
	if(x==?20'b111?????111????????0) z |= 4'b1000; 
	if(x==?20'b1?1?1?1?1?1????????0) z |= 4'b1000; 
	if(x==?20'b111???1?1?1????????0) z |= 4'b1000; 
	if(x==?20'b?1?1???1?111???????0) z |= 4'b0100; 
	if(x==?20'b?111?????111???????0) z |= 4'b0100; 
	if(x==?20'b?1?1?1?1?1?1???????0) z |= 4'b0100; 
	if(x==?20'b?111?1???1?1???????0) z |= 4'b0100; 
	if(x==?20'b????1?1???1?111????0) z |= 4'b0010; 
	if(x==?20'b????111?????111????0) z |= 4'b0010; 
	if(x==?20'b????1?1?1?1?1?1????0) z |= 4'b0010; 
	if(x==?20'b????111?1???1?1????0) z |= 4'b0010; 
	if(x==?20'b?????1?1?1???111???0) z |= 4'b0001; 
	if(x==?20'b?????111?????111???0) z |= 4'b0001; 
	if(x==?20'b?????1?1?1?1?1?1???0) z |= 4'b0001; 
	if(x==?20'b?????111???1?1?1???0) z |= 4'b0001; 
	if(x==?20'b??1??1??111?????000?) z |= 4'b1000; 
	if(x==?20'b?1??1?1??11?????000?) z |= 4'b1000; 
	if(x==?20'b??1??11?1?1?????000?) z |= 4'b1000; 
	if(x==?20'b?1????1??111????000?) z |= 4'b0100; 
	if(x==?20'b?1???11??1?1????000?) z |= 4'b0100; 
	if(x==?20'b??1??1?1?11?????000?) z |= 4'b0100; 
	if(x==?20'b????1?1??11???1?000?) z |= 4'b0010; 
	if(x==?20'b????111??1????1?000?) z |= 4'b0010; 
	if(x==?20'b?????11?1?1??1??000?) z |= 4'b0010; 
	if(x==?20'b?????11??1?1??1?000?) z |= 4'b0001; 
	if(x==?20'b?????1?1?11??1??000?) z |= 4'b0001; 
	if(x==?20'b?????111??1??1??000?) z |= 4'b0001; 
	if(x==?20'b??1??11?111?????0?0?) z |= 4'b1000; 
	if(x==?20'b?1???11??111????0?0?) z |= 4'b0100; 
	if(x==?20'b????111??11???1?0?0?) z |= 4'b0010; 
	if(x==?20'b?????111?11??1??0?0?) z |= 4'b0001; 
	if(x==?20'b?1??111??11?????00??) z |= 4'b1000; 
	if(x==?20'b??1??111?11?????00??) z |= 4'b0100; 
	if(x==?20'b?????11?111??1??00??) z |= 4'b0010; 
	if(x==?20'b?????11??111??1?00??) z |= 4'b0001; 
	if(x==?20'b?11?11??1????????00?) z |= 4'b1000; 
	if(x==?20'b?11???11???1?????00?) z |= 4'b0100; 
	if(x==?20'b????1???11???11??00?) z |= 4'b0010; 
	if(x==?20'b???????1??11?11??00?) z |= 4'b0001; 
	if(x==?20'b?11?11??11????????0?) z |= 4'b1000; 
	if(x==?20'b?11?111?1?????????0?) z |= 4'b1000; 
	if(x==?20'b?11???11??11??????0?) z |= 4'b0100; 
	if(x==?20'b?11??111???1??????0?) z |= 4'b0100; 
	if(x==?20'b????1???111??11???0?) z |= 4'b0010; 
	if(x==?20'b????11??11???11???0?) z |= 4'b0010; 
	if(x==?20'b???????1?111?11???0?) z |= 4'b0001; 
	if(x==?20'b??????11??11?11???0?) z |= 4'b0001; 
	if(x==?20'b?11?1???1?1?????0??0) z |= 4'b1000; 
	if(x==?20'b?11????1?1?1????0??0) z |= 4'b0100; 
	if(x==?20'b????1?1?1????11?0??0) z |= 4'b0010; 
	if(x==?20'b?????1?1???1?11?0??0) z |= 4'b0001; 
	if(x==?20'b11??11??????????000?) z |= 4'b1000; 
	if(x==?20'b??11??11????????000?) z |= 4'b0100; 
	if(x==?20'b????????11??11??000?) z |= 4'b0010; 
	if(x==?20'b??????????11??11000?) z |= 4'b0001; 
	if(x==?20'b11??11????1??????00?) z |= 4'b1000; 
	if(x==?20'b1???11??11???????00?) z |= 4'b1000; 
	if(x==?20'b11???1??11???????00?) z |= 4'b1000; 
	if(x==?20'b1?1?11???1???????00?) z |= 4'b1000; 
	if(x==?20'b111??1???1???????00?) z |= 4'b1000; 
	if(x==?20'b1???111?1????????00?) z |= 4'b1000; 
	if(x==?20'b11???11?1????????00?) z |= 4'b1000; 
	if(x==?20'b1?1?111??????????00?) z |= 4'b1000; 
	if(x==?20'b111??11??????????00?) z |= 4'b1000; 
	if(x==?20'b11??11???1??????0?0?) z |= 4'b1000; 
	if(x==?20'b11??111?????????0?0?) z |= 4'b1000; 
	if(x==?20'b???1??11??11?????00?) z |= 4'b0100; 
	if(x==?20'b??11??1???11?????00?) z |= 4'b0100; 
	if(x==?20'b???1?111???1?????00?) z |= 4'b0100; 
	if(x==?20'b??11?11????1?????00?) z |= 4'b0100; 
	if(x==?20'b?1?1??11??1??????00?) z |= 4'b0100; 
	if(x==?20'b?111??1???1??????00?) z |= 4'b0100; 
	if(x==?20'b??11??11?1???????00?) z |= 4'b0100; 
	if(x==?20'b?1?1?111?????????00?) z |= 4'b0100; 
	if(x==?20'b?111?11??????????00?) z |= 4'b0100; 
	if(x==?20'b??11??11??1?????0?0?) z |= 4'b0100; 
	if(x==?20'b??11?111????????0?0?) z |= 4'b0100; 
	if(x==?20'b?????????11?111??00?) z |= 4'b0010; 
	if(x==?20'b?????1???1??111??00?) z |= 4'b0010; 
	if(x==?20'b????????111?1?1??00?) z |= 4'b0010; 
	if(x==?20'b?????1??11??1?1??00?) z |= 4'b0010; 
	if(x==?20'b????1????11?11???00?) z |= 4'b0010; 
	if(x==?20'b??????1?11??11???00?) z |= 4'b0010; 
	if(x==?20'b????11???1??11???00?) z |= 4'b0010; 
	if(x==?20'b????1???111?1????00?) z |= 4'b0010; 
	if(x==?20'b????11??11??1????00?) z |= 4'b0010; 
	if(x==?20'b????????111?11??0?0?) z |= 4'b0010; 
	if(x==?20'b?????1??11??11??0?0?) z |= 4'b0010; 
	if(x==?20'b?????????11??111?00?) z |= 4'b0001; 
	if(x==?20'b??????1???1??111?00?) z |= 4'b0001; 
	if(x==?20'b?????1????11??11?00?) z |= 4'b0001; 
	if(x==?20'b???????1?11???11?00?) z |= 4'b0001; 
	if(x==?20'b??????11??1???11?00?) z |= 4'b0001; 
	if(x==?20'b?????????111?1?1?00?) z |= 4'b0001; 
	if(x==?20'b??????1???11?1?1?00?) z |= 4'b0001; 
	if(x==?20'b???????1?111???1?00?) z |= 4'b0001; 
	if(x==?20'b??????11??11???1?00?) z |= 4'b0001; 
	if(x==?20'b?????????111??110?0?) z |= 4'b0001; 
	if(x==?20'b??????1???11??110?0?) z |= 4'b0001; 
	if(x==?20'b11??11???11???????0?) z |= 4'b1000; 
	if(x==?20'b11??111???1???????0?) z |= 4'b1000; 
	if(x==?20'b1???111?11????????0?) z |= 4'b1000; 
	if(x==?20'b11???11?11????????0?) z |= 4'b1000; 
	if(x==?20'b1?1?111??1????????0?) z |= 4'b1000; 
	if(x==?20'b111??11??1????????0?) z |= 4'b1000; 
	if(x==?20'b???1?111??11??????0?) z |= 4'b0100; 
	if(x==?20'b??11?11???11??????0?) z |= 4'b0100; 
	if(x==?20'b??11??11?11???????0?) z |= 4'b0100; 
	if(x==?20'b?1?1?111??1???????0?) z |= 4'b0100; 
	if(x==?20'b?111?11???1???????0?) z |= 4'b0100; 
	if(x==?20'b??11?111?1????????0?) z |= 4'b0100; 
	if(x==?20'b?????1???11?111???0?) z |= 4'b0010; 
	if(x==?20'b?????1??111?1?1???0?) z |= 4'b0010; 
	if(x==?20'b??????1?111?11????0?) z |= 4'b0010; 
	if(x==?20'b????11???11?11????0?) z |= 4'b0010; 
	if(x==?20'b?????11?11??11????0?) z |= 4'b0010; 
	if(x==?20'b????11??111?1?????0?) z |= 4'b0010; 
	if(x==?20'b??????1??11??111??0?) z |= 4'b0001; 
	if(x==?20'b?????1???111??11??0?) z |= 4'b0001; 
	if(x==?20'b?????11???11??11??0?) z |= 4'b0001; 
	if(x==?20'b??????11?11???11??0?) z |= 4'b0001; 
	if(x==?20'b??????1??111?1?1??0?) z |= 4'b0001; 
	if(x==?20'b??????11?111???1??0?) z |= 4'b0001; 
	if(x==?20'b1???1???1?1?????00?0) z |= 4'b1000; 
	if(x==?20'b11??????1?1?????00?0) z |= 4'b1000; 
	if(x==?20'b1?1?1?????1?????00?0) z |= 4'b1000; 
	if(x==?20'b111???????1?????00?0) z |= 4'b1000; 
	if(x==?20'b1?1?????11??????00?0) z |= 4'b1000; 
	if(x==?20'b1?1???1?1???????00?0) z |= 4'b1000; 
	if(x==?20'b?1?1??????11????00?0) z |= 4'b0100; 
	if(x==?20'b???1???1?1?1????00?0) z |= 4'b0100; 
	if(x==?20'b??11?????1?1????00?0) z |= 4'b0100; 
	if(x==?20'b?1?1?1?????1????00?0) z |= 4'b0100; 
	if(x==?20'b?1?1???1?1??????00?0) z |= 4'b0100; 
	if(x==?20'b?111?????1??????00?0) z |= 4'b0100; 
	if(x==?20'b??????1?????111?00?0) z |= 4'b0010; 
	if(x==?20'b????1?????1?1?1?00?0) z |= 4'b0010; 
	if(x==?20'b??????1?1???1?1?00?0) z |= 4'b0010; 
	if(x==?20'b????11??????1?1?00?0) z |= 4'b0010; 
	if(x==?20'b????1?1?????11??00?0) z |= 4'b0010; 
	if(x==?20'b????1?1?1???1???00?0) z |= 4'b0010; 
	if(x==?20'b?????1???????11100?0) z |= 4'b0001; 
	if(x==?20'b?????1?1??????1100?0) z |= 4'b0001; 
	if(x==?20'b?????1?????1?1?100?0) z |= 4'b0001; 
	if(x==?20'b???????1?1???1?100?0) z |= 4'b0001; 
	if(x==?20'b??????11?????1?100?0) z |= 4'b0001; 
	if(x==?20'b?????1?1???1???100?0) z |= 4'b0001; 
	if(x==?20'b1?1?????111??????0?0) z |= 4'b1000; 
	if(x==?20'b1?1???1?1?1??????0?0) z |= 4'b1000; 
	if(x==?20'b1???1???111?????0??0) z |= 4'b1000; 
	if(x==?20'b11??????111?????0??0) z |= 4'b1000; 
	if(x==?20'b1?1?1????11?????0??0) z |= 4'b1000; 
	if(x==?20'b111??????11?????0??0) z |= 4'b1000; 
	if(x==?20'b1???1?1?1?1?????0??0) z |= 4'b1000; 
	if(x==?20'b11????1?1?1?????0??0) z |= 4'b1000; 
	if(x==?20'b1?1?1?1???1?????0??0) z |= 4'b1000; 
	if(x==?20'b111???1???1?????0??0) z |= 4'b1000; 
	if(x==?20'b1?1???1?11??????0??0) z |= 4'b1000; 
	if(x==?20'b?1?1?????111?????0?0) z |= 4'b0100; 
	if(x==?20'b?1?1?1???1?1?????0?0) z |= 4'b0100; 
	if(x==?20'b???1???1?111????0??0) z |= 4'b0100; 
	if(x==?20'b??11?????111????0??0) z |= 4'b0100; 
	if(x==?20'b?1?1?1????11????0??0) z |= 4'b0100; 
	if(x==?20'b???1?1?1?1?1????0??0) z |= 4'b0100; 
	if(x==?20'b??11?1???1?1????0??0) z |= 4'b0100; 
	if(x==?20'b?1?1???1?11?????0??0) z |= 4'b0100; 
	if(x==?20'b?111?????11?????0??0) z |= 4'b0100; 
	if(x==?20'b?1?1?1?1?1??????0??0) z |= 4'b0100; 
	if(x==?20'b?111?1???1??????0??0) z |= 4'b0100; 
	if(x==?20'b????1?1???1?1?1??0?0) z |= 4'b0010; 
	if(x==?20'b????111?????1?1??0?0) z |= 4'b0010; 
	if(x==?20'b??????1???1?111?0??0) z |= 4'b0010; 
	if(x==?20'b?????11?????111?0??0) z |= 4'b0010; 
	if(x==?20'b??????1?1?1?1?1?0??0) z |= 4'b0010; 
	if(x==?20'b????11????1?1?1?0??0) z |= 4'b0010; 
	if(x==?20'b?????11?1???1?1?0??0) z |= 4'b0010; 
	if(x==?20'b????1?1???1?11??0??0) z |= 4'b0010; 
	if(x==?20'b????111?????11??0??0) z |= 4'b0010; 
	if(x==?20'b????1?1?1?1?1???0??0) z |= 4'b0010; 
	if(x==?20'b????111?1???1???0??0) z |= 4'b0010; 
	if(x==?20'b?????1?1?1???1?1?0?0) z |= 4'b0001; 
	if(x==?20'b?????111?????1?1?0?0) z |= 4'b0001; 
	if(x==?20'b?????1???1???1110??0) z |= 4'b0001; 
	if(x==?20'b?????11??????1110??0) z |= 4'b0001; 
	if(x==?20'b?????1?1?1????110??0) z |= 4'b0001; 
	if(x==?20'b?????111??????110??0) z |= 4'b0001; 
	if(x==?20'b?????1???1?1?1?10??0) z |= 4'b0001; 
	if(x==?20'b?????11????1?1?10??0) z |= 4'b0001; 
	if(x==?20'b??????11?1???1?10??0) z |= 4'b0001; 
	if(x==?20'b?????1?1?1?1???10??0) z |= 4'b0001; 
	if(x==?20'b?????111???1???10??0) z |= 4'b0001; 
	if(x==?20'b1?1???1?111????????0) z |= 4'b1000; 
	if(x==?20'b?1?1?1???111???????0) z |= 4'b0100; 
	if(x==?20'b????111???1?1?1????0) z |= 4'b0010; 
	if(x==?20'b?????111?1???1?1???0) z |= 4'b0001; 
	if(x==?20'b?1??11??1???????000?) z |= 4'b1000; 
	if(x==?20'b?11?11??????????000?) z |= 4'b1000; 
	if(x==?20'b??1???11???1????000?) z |= 4'b0100; 
	if(x==?20'b?11???11????????000?) z |= 4'b0100; 
	if(x==?20'b????????11???11?000?) z |= 4'b0010; 
	if(x==?20'b????1???11???1??000?) z |= 4'b0010; 
	if(x==?20'b??????????11?11?000?) z |= 4'b0001; 
	if(x==?20'b???????1??11??1?000?) z |= 4'b0001; 
	if(x==?20'b?1??11??1?1??????00?) z |= 4'b1000; 
	if(x==?20'b?11?11????1??????00?) z |= 4'b1000; 
	if(x==?20'b??1?11??11???????00?) z |= 4'b1000; 
	if(x==?20'b?11??1??11???????00?) z |= 4'b1000; 
	if(x==?20'b??1?111?1????????00?) z |= 4'b1000; 
	if(x==?20'b?11??11?1????????00?) z |= 4'b1000; 
	if(x==?20'b?1??11??11??????0?0?) z |= 4'b1000; 
	if(x==?20'b?11?11???1??????0?0?) z |= 4'b1000; 
	if(x==?20'b?1??111?1???????0?0?) z |= 4'b1000; 
	if(x==?20'b?11?111?????????0?0?) z |= 4'b1000; 
	if(x==?20'b?1????11??11?????00?) z |= 4'b0100; 
	if(x==?20'b?11???1???11?????00?) z |= 4'b0100; 
	if(x==?20'b??1???11?1?1?????00?) z |= 4'b0100; 
	if(x==?20'b?1???111???1?????00?) z |= 4'b0100; 
	if(x==?20'b?11??11????1?????00?) z |= 4'b0100; 
	if(x==?20'b?11???11?1???????00?) z |= 4'b0100; 
	if(x==?20'b??1???11??11????0?0?) z |= 4'b0100; 
	if(x==?20'b??1??111???1????0?0?) z |= 4'b0100; 
	if(x==?20'b?11???11??1?????0?0?) z |= 4'b0100; 
	if(x==?20'b?11??111????????0?0?) z |= 4'b0100; 
	if(x==?20'b????1????11??11??00?) z |= 4'b0010; 
	if(x==?20'b??????1?11???11??00?) z |= 4'b0010; 
	if(x==?20'b????11???1???11??00?) z |= 4'b0010; 
	if(x==?20'b????1???111???1??00?) z |= 4'b0010; 
	if(x==?20'b????11??11????1??00?) z |= 4'b0010; 
	if(x==?20'b????1?1?11???1???00?) z |= 4'b0010; 
	if(x==?20'b????????111??11?0?0?) z |= 4'b0010; 
	if(x==?20'b?????1??11???11?0?0?) z |= 4'b0010; 
	if(x==?20'b????1???111??1??0?0?) z |= 4'b0010; 
	if(x==?20'b????11??11???1??0?0?) z |= 4'b0010; 
	if(x==?20'b?????1????11?11??00?) z |= 4'b0001; 
	if(x==?20'b???????1?11??11??00?) z |= 4'b0001; 
	if(x==?20'b??????11??1??11??00?) z |= 4'b0001; 
	if(x==?20'b?????1?1??11??1??00?) z |= 4'b0001; 
	if(x==?20'b???????1?111?1???00?) z |= 4'b0001; 
	if(x==?20'b??????11??11?1???00?) z |= 4'b0001; 
	if(x==?20'b?????????111?11?0?0?) z |= 4'b0001; 
	if(x==?20'b??????1???11?11?0?0?) z |= 4'b0001; 
	if(x==?20'b???????1?111??1?0?0?) z |= 4'b0001; 
	if(x==?20'b??????11??11??1?0?0?) z |= 4'b0001; 
	if(x==?20'b?1??11??111???????0?) z |= 4'b1000; 
	if(x==?20'b?11?11???11???????0?) z |= 4'b1000; 
	if(x==?20'b?1??111?1?1???????0?) z |= 4'b1000; 
	if(x==?20'b?11?111???1???????0?) z |= 4'b1000; 
	if(x==?20'b??1?111?11????????0?) z |= 4'b1000; 
	if(x==?20'b?11??11?11????????0?) z |= 4'b1000; 
	if(x==?20'b??1???11?111??????0?) z |= 4'b0100; 
	if(x==?20'b?1???111??11??????0?) z |= 4'b0100; 
	if(x==?20'b?11??11???11??????0?) z |= 4'b0100; 
	if(x==?20'b??1??111?1?1??????0?) z |= 4'b0100; 
	if(x==?20'b?11???11?11???????0?) z |= 4'b0100; 
	if(x==?20'b?11??111?1????????0?) z |= 4'b0100; 
	if(x==?20'b??????1?111??11???0?) z |= 4'b0010; 
	if(x==?20'b????11???11??11???0?) z |= 4'b0010; 
	if(x==?20'b?????11?11???11???0?) z |= 4'b0010; 
	if(x==?20'b????11??111???1???0?) z |= 4'b0010; 
	if(x==?20'b????1?1?111??1????0?) z |= 4'b0010; 
	if(x==?20'b????111?11???1????0?) z |= 4'b0010; 
	if(x==?20'b?????1???111?11???0?) z |= 4'b0001; 
	if(x==?20'b?????11???11?11???0?) z |= 4'b0001; 
	if(x==?20'b??????11?11??11???0?) z |= 4'b0001; 
	if(x==?20'b?????1?1?111??1???0?) z |= 4'b0001; 
	if(x==?20'b?????111??11??1???0?) z |= 4'b0001; 
	if(x==?20'b??????11?111?1????0?) z |= 4'b0001; 
	if(x==?20'b??1?1???1?1?????00?0) z |= 4'b1000; 
	if(x==?20'b?11?????1?1?????00?0) z |= 4'b1000; 
	if(x==?20'b?1?????1?1?1????00?0) z |= 4'b0100; 
	if(x==?20'b?11??????1?1????00?0) z |= 4'b0100; 
	if(x==?20'b????1?1??????11?00?0) z |= 4'b0010; 
	if(x==?20'b????1?1?1?????1?00?0) z |= 4'b0010; 
	if(x==?20'b?????1?1?????11?00?0) z |= 4'b0001; 
	if(x==?20'b?????1?1???1?1??00?0) z |= 4'b0001; 
	if(x==?20'b??1?1???111?????0??0) z |= 4'b1000; 
	if(x==?20'b?11?????111?????0??0) z |= 4'b1000; 
	if(x==?20'b??1?1?1?1?1?????0??0) z |= 4'b1000; 
	if(x==?20'b?11???1?1?1?????0??0) z |= 4'b1000; 
	if(x==?20'b?1?????1?111????0??0) z |= 4'b0100; 
	if(x==?20'b?11??????111????0??0) z |= 4'b0100; 
	if(x==?20'b?1???1?1?1?1????0??0) z |= 4'b0100; 
	if(x==?20'b?11??1???1?1????0??0) z |= 4'b0100; 
	if(x==?20'b????1?1???1??11?0??0) z |= 4'b0010; 
	if(x==?20'b????111??????11?0??0) z |= 4'b0010; 
	if(x==?20'b????1?1?1?1???1?0??0) z |= 4'b0010; 
	if(x==?20'b????111?1?????1?0??0) z |= 4'b0010; 
	if(x==?20'b?????1?1?1???11?0??0) z |= 4'b0001; 
	if(x==?20'b?????111?????11?0??0) z |= 4'b0001; 
	if(x==?20'b?????1?1?1?1?1??0??0) z |= 4'b0001; 
	if(x==?20'b?????111???1?1??0??0) z |= 4'b0001; 
	if(x==?20'b1???11???1??????000?) z |= 4'b1000; 
	if(x==?20'b11???1???1??????000?) z |= 4'b1000; 
	if(x==?20'b1???111?????????000?) z |= 4'b1000; 
	if(x==?20'b11???11?????????000?) z |= 4'b1000; 
	if(x==?20'b???1??11??1?????000?) z |= 4'b0100; 
	if(x==?20'b??11??1???1?????000?) z |= 4'b0100; 
	if(x==?20'b???1?111????????000?) z |= 4'b0100; 
	if(x==?20'b??11?11?????????000?) z |= 4'b0100; 
	if(x==?20'b?????????11?11??000?) z |= 4'b0010; 
	if(x==?20'b?????1???1??11??000?) z |= 4'b0010; 
	if(x==?20'b????????111?1???000?) z |= 4'b0010; 
	if(x==?20'b?????1??11??1???000?) z |= 4'b0010; 
	if(x==?20'b?????????11???11000?) z |= 4'b0001; 
	if(x==?20'b??????1???1???11000?) z |= 4'b0001; 
	if(x==?20'b?????????111???1000?) z |= 4'b0001; 
	if(x==?20'b??????1???11???1000?) z |= 4'b0001; 
	if(x==?20'b1???11???11??????00?) z |= 4'b1000; 
	if(x==?20'b11???1???11??????00?) z |= 4'b1000; 
	if(x==?20'b1???111???1??????00?) z |= 4'b1000; 
	if(x==?20'b11???11???1??????00?) z |= 4'b1000; 
	if(x==?20'b1????11?11???????00?) z |= 4'b1000; 
	if(x==?20'b1?1??11??1???????00?) z |= 4'b1000; 
	if(x==?20'b1???111??1??????0?0?) z |= 4'b1000; 
	if(x==?20'b11???11??1??????0?0?) z |= 4'b1000; 
	if(x==?20'b???1?11???11?????00?) z |= 4'b0100; 
	if(x==?20'b???1??11?11??????00?) z |= 4'b0100; 
	if(x==?20'b??11??1??11??????00?) z |= 4'b0100; 
	if(x==?20'b?1?1?11???1??????00?) z |= 4'b0100; 
	if(x==?20'b???1?111?1???????00?) z |= 4'b0100; 
	if(x==?20'b??11?11??1???????00?) z |= 4'b0100; 
	if(x==?20'b???1?111??1?????0?0?) z |= 4'b0100; 
	if(x==?20'b??11?11???1?????0?0?) z |= 4'b0100; 
	if(x==?20'b?????1???11?1?1??00?) z |= 4'b0010; 
	if(x==?20'b??????1??11?11???00?) z |= 4'b0010; 
	if(x==?20'b?????11??1??11???00?) z |= 4'b0010; 
	if(x==?20'b??????1?111?1????00?) z |= 4'b0010; 
	if(x==?20'b????11???11?1????00?) z |= 4'b0010; 
	if(x==?20'b?????11?11??1????00?) z |= 4'b0010; 
	if(x==?20'b?????1???11?11??0?0?) z |= 4'b0010; 
	if(x==?20'b?????1??111?1???0?0?) z |= 4'b0010; 
	if(x==?20'b?????1???11???11?00?) z |= 4'b0001; 
	if(x==?20'b?????11???1???11?00?) z |= 4'b0001; 
	if(x==?20'b??????1??11??1?1?00?) z |= 4'b0001; 
	if(x==?20'b?????1???111???1?00?) z |= 4'b0001; 
	if(x==?20'b?????11???11???1?00?) z |= 4'b0001; 
	if(x==?20'b??????11?11????1?00?) z |= 4'b0001; 
	if(x==?20'b??????1??11???110?0?) z |= 4'b0001; 
	if(x==?20'b??????1??111???10?0?) z |= 4'b0001; 
	if(x==?20'b1???111??11???????0?) z |= 4'b1000; 
	if(x==?20'b11???11??11???????0?) z |= 4'b1000; 
	if(x==?20'b???1?111?11???????0?) z |= 4'b0100; 
	if(x==?20'b??11?11??11???????0?) z |= 4'b0100; 
	if(x==?20'b?????11??11?11????0?) z |= 4'b0010; 
	if(x==?20'b?????11?111?1?????0?) z |= 4'b0010; 
	if(x==?20'b?????11??11???11??0?) z |= 4'b0001; 
	if(x==?20'b?????11??111???1??0?) z |= 4'b0001; 
	if(x==?20'b1???????111?????00?0) z |= 4'b1000; 
	if(x==?20'b1?1??????11?????00?0) z |= 4'b1000; 
	if(x==?20'b1?????1?1?1?????00?0) z |= 4'b1000; 
	if(x==?20'b1?1???1???1?????00?0) z |= 4'b1000; 
	if(x==?20'b???1?????111????00?0) z |= 4'b0100; 
	if(x==?20'b???1?1???1?1????00?0) z |= 4'b0100; 
	if(x==?20'b?1?1?????11?????00?0) z |= 4'b0100; 
	if(x==?20'b?1?1?1???1??????00?0) z |= 4'b0100; 
	if(x==?20'b??????1???1?1?1?00?0) z |= 4'b0010; 
	if(x==?20'b?????11?????1?1?00?0) z |= 4'b0010; 
	if(x==?20'b????1?1???1?1???00?0) z |= 4'b0010; 
	if(x==?20'b????111?????1???00?0) z |= 4'b0010; 
	if(x==?20'b?????1???1???1?100?0) z |= 4'b0001; 
	if(x==?20'b?????11??????1?100?0) z |= 4'b0001; 
	if(x==?20'b?????1?1?1?????100?0) z |= 4'b0001; 
	if(x==?20'b?????111???????100?0) z |= 4'b0001; 
	if(x==?20'b1?????1?111?????0??0) z |= 4'b1000; 
	if(x==?20'b1?1???1??11?????0??0) z |= 4'b1000; 
	if(x==?20'b???1?1???111????0??0) z |= 4'b0100; 
	if(x==?20'b?1?1?1???11?????0??0) z |= 4'b0100; 
	if(x==?20'b?????11???1?1?1?0??0) z |= 4'b0010; 
	if(x==?20'b????111???1?1???0??0) z |= 4'b0010; 
	if(x==?20'b?????11??1???1?10??0) z |= 4'b0001; 
	if(x==?20'b?????111?1?????10??0) z |= 4'b0001; 
	if(x==?20'b11??1???1????????0?0) z |= 4'b1000; 
	if(x==?20'b111?1????????????0?0) z |= 4'b1000; 
	if(x==?20'b??11???1???1?????0?0) z |= 4'b0100; 
	if(x==?20'b?111???1?????????0?0) z |= 4'b0100; 
	if(x==?20'b????????1???111??0?0) z |= 4'b0010; 
	if(x==?20'b????1???1???11???0?0) z |= 4'b0010; 
	if(x==?20'b???????????1?111?0?0) z |= 4'b0001; 
	if(x==?20'b???????1???1??11?0?0) z |= 4'b0001; 
	if(x==?20'b11??1???11?????????0) z |= 4'b1000; 
	if(x==?20'b111?1????1?????????0) z |= 4'b1000; 
	if(x==?20'b11??1?1?1??????????0) z |= 4'b1000; 
	if(x==?20'b111?1?1????????????0) z |= 4'b1000; 
	if(x==?20'b??11???1??11???????0) z |= 4'b0100; 
	if(x==?20'b??11?1?1???1???????0) z |= 4'b0100; 
	if(x==?20'b?111???1??1????????0) z |= 4'b0100; 
	if(x==?20'b?111?1?1???????????0) z |= 4'b0100; 
	if(x==?20'b????????1?1?111????0) z |= 4'b0010; 
	if(x==?20'b?????1??1???111????0) z |= 4'b0010; 
	if(x==?20'b????1???1?1?11?????0) z |= 4'b0010; 
	if(x==?20'b????11??1???11?????0) z |= 4'b0010; 
	if(x==?20'b?????????1?1?111???0) z |= 4'b0001; 
	if(x==?20'b??????1????1?111???0) z |= 4'b0001; 
	if(x==?20'b???????1?1?1??11???0) z |= 4'b0001; 
	if(x==?20'b??????11???1??11???0) z |= 4'b0001; 
	if(x==?20'b?1??11????1?????000?) z |= 4'b1000; 
	if(x==?20'b?1???1??11??????000?) z |= 4'b1000; 
	if(x==?20'b??1?11???1??????000?) z |= 4'b1000; 
	if(x==?20'b?11??1???1??????000?) z |= 4'b1000; 
	if(x==?20'b????111?1???????000?) z |= 4'b1000; 
	if(x==?20'b?1???11?1???????000?) z |= 4'b1000; 
	if(x==?20'b??1?111?????????000?) z |= 4'b1000; 
	if(x==?20'b??1???1???11????000?) z |= 4'b0100; 
	if(x==?20'b?????111???1????000?) z |= 4'b0100; 
	if(x==?20'b??1??11????1????000?) z |= 4'b0100; 
	if(x==?20'b?1????11??1?????000?) z |= 4'b0100; 
	if(x==?20'b?11???1???1?????000?) z |= 4'b0100; 
	if(x==?20'b??1???11?1??????000?) z |= 4'b0100; 
	if(x==?20'b?1???111????????000?) z |= 4'b0100; 
	if(x==?20'b?????1???1???11?000?) z |= 4'b0010; 
	if(x==?20'b????????111???1?000?) z |= 4'b0010; 
	if(x==?20'b?????1??11????1?000?) z |= 4'b0010; 
	if(x==?20'b????1????11??1??000?) z |= 4'b0010; 
	if(x==?20'b??????1?11???1??000?) z |= 4'b0010; 
	if(x==?20'b????11???1???1??000?) z |= 4'b0010; 
	if(x==?20'b????1???111?????000?) z |= 4'b0010; 
	if(x==?20'b??????1???1??11?000?) z |= 4'b0001; 
	if(x==?20'b?????1????11??1?000?) z |= 4'b0001; 
	if(x==?20'b???????1?11???1?000?) z |= 4'b0001; 
	if(x==?20'b??????11??1???1?000?) z |= 4'b0001; 
	if(x==?20'b?????????111?1??000?) z |= 4'b0001; 
	if(x==?20'b??????1???11?1??000?) z |= 4'b0001; 
	if(x==?20'b???????1?111????000?) z |= 4'b0001; 
	if(x==?20'b????11??111??????00?) z |= 4'b1000; 
	if(x==?20'b?1???1??111??????00?) z |= 4'b1000; 
	if(x==?20'b??1?11???11??????00?) z |= 4'b1000; 
	if(x==?20'b?11??1???11??????00?) z |= 4'b1000; 
	if(x==?20'b????111?1?1??????00?) z |= 4'b1000; 
	if(x==?20'b?1???11?1?1??????00?) z |= 4'b1000; 
	if(x==?20'b??1?111???1??????00?) z |= 4'b1000; 
	if(x==?20'b?11??11???1??????00?) z |= 4'b1000; 
	if(x==?20'b??1??11?11???????00?) z |= 4'b1000; 
	if(x==?20'b?1??11???11?????0?0?) z |= 4'b1000; 
	if(x==?20'b?1??111???1?????0?0?) z |= 4'b1000; 
	if(x==?20'b????111?11??????0?0?) z |= 4'b1000; 
	if(x==?20'b?1???11?11??????0?0?) z |= 4'b1000; 
	if(x==?20'b??1?111??1??????0?0?) z |= 4'b1000; 
	if(x==?20'b?11??11??1??????0?0?) z |= 4'b1000; 
	if(x==?20'b??????11?111?????00?) z |= 4'b0100; 
	if(x==?20'b??1???1??111?????00?) z |= 4'b0100; 
	if(x==?20'b?1???11???11?????00?) z |= 4'b0100; 
	if(x==?20'b?????111?1?1?????00?) z |= 4'b0100; 
	if(x==?20'b??1??11??1?1?????00?) z |= 4'b0100; 
	if(x==?20'b?1????11?11??????00?) z |= 4'b0100; 
	if(x==?20'b?11???1??11??????00?) z |= 4'b0100; 
	if(x==?20'b?1???111?1???????00?) z |= 4'b0100; 
	if(x==?20'b?11??11??1???????00?) z |= 4'b0100; 
	if(x==?20'b?????111??11????0?0?) z |= 4'b0100; 
	if(x==?20'b??1??11???11????0?0?) z |= 4'b0100; 
	if(x==?20'b??1???11?11?????0?0?) z |= 4'b0100; 
	if(x==?20'b?1???111??1?????0?0?) z |= 4'b0100; 
	if(x==?20'b?11??11???1?????0?0?) z |= 4'b0100; 
	if(x==?20'b??1??111?1??????0?0?) z |= 4'b0100; 
	if(x==?20'b??????1??11??11??00?) z |= 4'b0010; 
	if(x==?20'b?????11??1???11??00?) z |= 4'b0010; 
	if(x==?20'b??????1?111???1??00?) z |= 4'b0010; 
	if(x==?20'b????11???11???1??00?) z |= 4'b0010; 
	if(x==?20'b?????11?11????1??00?) z |= 4'b0010; 
	if(x==?20'b????1?1??11??1???00?) z |= 4'b0010; 
	if(x==?20'b????111??1???1???00?) z |= 4'b0010; 
	if(x==?20'b????1?1?111??????00?) z |= 4'b0010; 
	if(x==?20'b????111?11???????00?) z |= 4'b0010; 
	if(x==?20'b?????1???11??11?0?0?) z |= 4'b0010; 
	if(x==?20'b?????1??111???1?0?0?) z |= 4'b0010; 
	if(x==?20'b??????1?111??1??0?0?) z |= 4'b0010; 
	if(x==?20'b????11???11??1??0?0?) z |= 4'b0010; 
	if(x==?20'b?????11?11???1??0?0?) z |= 4'b0010; 
	if(x==?20'b????11??111?????0?0?) z |= 4'b0010; 
	if(x==?20'b?????1???11??11??00?) z |= 4'b0001; 
	if(x==?20'b?????11???1??11??00?) z |= 4'b0001; 
	if(x==?20'b?????1?1?11???1??00?) z |= 4'b0001; 
	if(x==?20'b?????111??1???1??00?) z |= 4'b0001; 
	if(x==?20'b?????1???111?1???00?) z |= 4'b0001; 
	if(x==?20'b?????11???11?1???00?) z |= 4'b0001; 
	if(x==?20'b??????11?11??1???00?) z |= 4'b0001; 
	if(x==?20'b?????1?1?111?????00?) z |= 4'b0001; 
	if(x==?20'b?????111??11?????00?) z |= 4'b0001; 
	if(x==?20'b??????1??11??11?0?0?) z |= 4'b0001; 
	if(x==?20'b?????1???111??1?0?0?) z |= 4'b0001; 
	if(x==?20'b?????11???11??1?0?0?) z |= 4'b0001; 
	if(x==?20'b??????11?11???1?0?0?) z |= 4'b0001; 
	if(x==?20'b??????1??111?1??0?0?) z |= 4'b0001; 
	if(x==?20'b??????11?111????0?0?) z |= 4'b0001; 
	if(x==?20'b?1???11?111???????0?) z |= 4'b1000; 
	if(x==?20'b??1?111??11???????0?) z |= 4'b1000; 
	if(x==?20'b??1??11??111??????0?) z |= 4'b0100; 
	if(x==?20'b?1???111?11???????0?) z |= 4'b0100; 
	if(x==?20'b?????11?111???1???0?) z |= 4'b0010; 
	if(x==?20'b????111??11??1????0?) z |= 4'b0010; 
	if(x==?20'b?????111?11???1???0?) z |= 4'b0001; 
	if(x==?20'b?????11??111?1????0?) z |= 4'b0001; 
	if(x==?20'b??1?????111?????00?0) z |= 4'b1000; 
	if(x==?20'b??1???1?1?1?????00?0) z |= 4'b1000; 
	if(x==?20'b?1???????111????00?0) z |= 4'b0100; 
	if(x==?20'b?1???1???1?1????00?0) z |= 4'b0100; 
	if(x==?20'b????1?1???1???1?00?0) z |= 4'b0010; 
	if(x==?20'b????111???????1?00?0) z |= 4'b0010; 
	if(x==?20'b?????1?1?1???1??00?0) z |= 4'b0001; 
	if(x==?20'b?????111?????1??00?0) z |= 4'b0001; 
	if(x==?20'b??1???1?111?????0??0) z |= 4'b1000; 
	if(x==?20'b?1???1???111????0??0) z |= 4'b0100; 
	if(x==?20'b????111???1???1?0??0) z |= 4'b0010; 
	if(x==?20'b?????111?1???1??0??0) z |= 4'b0001; 
	if(x==?20'b?11?1???1????????0?0) z |= 4'b1000; 
	if(x==?20'b?11????1???1?????0?0) z |= 4'b0100; 
	if(x==?20'b????1???1????11??0?0) z |= 4'b0010; 
	if(x==?20'b???????1???1?11??0?0) z |= 4'b0001; 
	if(x==?20'b?11?1???11?????????0) z |= 4'b1000; 
	if(x==?20'b?11?1?1?1??????????0) z |= 4'b1000; 
	if(x==?20'b?11????1??11???????0) z |= 4'b0100; 
	if(x==?20'b?11??1?1???1???????0) z |= 4'b0100; 
	if(x==?20'b????1???1?1??11????0) z |= 4'b0010; 
	if(x==?20'b????11??1????11????0) z |= 4'b0010; 
	if(x==?20'b???????1?1?1?11????0) z |= 4'b0001; 
	if(x==?20'b??????11???1?11????0) z |= 4'b0001; 
	if(x==?20'b1????11??1??????000?) z |= 4'b1000; 
	if(x==?20'b???1?11???1?????000?) z |= 4'b0100; 
	if(x==?20'b?????1???11?1???000?) z |= 4'b0010; 
	if(x==?20'b??????1??11????1000?) z |= 4'b0001; 
	if(x==?20'b1????11??11??????00?) z |= 4'b1000; 
	if(x==?20'b???1?11??11??????00?) z |= 4'b0100; 
	if(x==?20'b?????11??11?1????00?) z |= 4'b0010; 
	if(x==?20'b?????11??11????1?00?) z |= 4'b0001; 
	if(x==?20'b1?1?????1???????0?00) z |= 4'b1000; 
	if(x==?20'b?1?1???????1????0?00) z |= 4'b0100; 
	if(x==?20'b????1???????1?1?0?00) z |= 4'b0010; 
	if(x==?20'b???????1?????1?10?00) z |= 4'b0001; 
	if(x==?20'b1?1?????1?1???????00) z |= 4'b1000; 
	if(x==?20'b11??1???????????00?0) z |= 4'b1000; 
	if(x==?20'b?1?1?????1?1??????00) z |= 4'b0100; 
	if(x==?20'b??11???1????????00?0) z |= 4'b0100; 
	if(x==?20'b????1?1?????1?1???00) z |= 4'b0010; 
	if(x==?20'b????????1???11??00?0) z |= 4'b0010; 
	if(x==?20'b?????1?1?????1?1??00) z |= 4'b0001; 
	if(x==?20'b???????????1??1100?0) z |= 4'b0001; 
	if(x==?20'b11??1?????1??????0?0) z |= 4'b1000; 
	if(x==?20'b1???1???11???????0?0) z |= 4'b1000; 
	if(x==?20'b11??????11???????0?0) z |= 4'b1000; 
	if(x==?20'b1?1?1????1???????0?0) z |= 4'b1000; 
	if(x==?20'b111??????1???????0?0) z |= 4'b1000; 
	if(x==?20'b1???1?1?1????????0?0) z |= 4'b1000; 
	if(x==?20'b11????1?1????????0?0) z |= 4'b1000; 
	if(x==?20'b1?1?1?1??????????0?0) z |= 4'b1000; 
	if(x==?20'b111???1??????????0?0) z |= 4'b1000; 
	if(x==?20'b11??1????1??????0??0) z |= 4'b1000; 
	if(x==?20'b1?1??1??1???????0??0) z |= 4'b1000; 
	if(x==?20'b11??1?1?????????0??0) z |= 4'b1000; 
	if(x==?20'b???1???1??11?????0?0) z |= 4'b0100; 
	if(x==?20'b??11??????11?????0?0) z |= 4'b0100; 
	if(x==?20'b???1?1?1???1?????0?0) z |= 4'b0100; 
	if(x==?20'b??11?1?????1?????0?0) z |= 4'b0100; 
	if(x==?20'b?1?1???1??1??????0?0) z |= 4'b0100; 
	if(x==?20'b?111??????1??????0?0) z |= 4'b0100; 
	if(x==?20'b??11???1?1???????0?0) z |= 4'b0100; 
	if(x==?20'b?1?1?1?1?????????0?0) z |= 4'b0100; 
	if(x==?20'b?111?1???????????0?0) z |= 4'b0100; 
	if(x==?20'b?1?1??1????1????0??0) z |= 4'b0100; 
	if(x==?20'b??11???1??1?????0??0) z |= 4'b0100; 
	if(x==?20'b??11?1?1????????0??0) z |= 4'b0100; 
	if(x==?20'b??????????1?111??0?0) z |= 4'b0010; 
	if(x==?20'b?????1??????111??0?0) z |= 4'b0010; 
	if(x==?20'b????????1?1?1?1??0?0) z |= 4'b0010; 
	if(x==?20'b?????1??1???1?1??0?0) z |= 4'b0010; 
	if(x==?20'b????1?????1?11???0?0) z |= 4'b0010; 
	if(x==?20'b??????1?1???11???0?0) z |= 4'b0010; 
	if(x==?20'b????11??????11???0?0) z |= 4'b0010; 
	if(x==?20'b????1???1?1?1????0?0) z |= 4'b0010; 
	if(x==?20'b????11??1???1????0?0) z |= 4'b0010; 
	if(x==?20'b????1????1??1?1?0??0) z |= 4'b0010; 
	if(x==?20'b????????1?1?11??0??0) z |= 4'b0010; 
	if(x==?20'b?????1??1???11??0??0) z |= 4'b0010; 
	if(x==?20'b?????????1???111?0?0) z |= 4'b0001; 
	if(x==?20'b??????1??????111?0?0) z |= 4'b0001; 
	if(x==?20'b?????1?????1??11?0?0) z |= 4'b0001; 
	if(x==?20'b???????1?1????11?0?0) z |= 4'b0001; 
	if(x==?20'b??????11??????11?0?0) z |= 4'b0001; 
	if(x==?20'b?????????1?1?1?1?0?0) z |= 4'b0001; 
	if(x==?20'b??????1????1?1?1?0?0) z |= 4'b0001; 
	if(x==?20'b???????1?1?1???1?0?0) z |= 4'b0001; 
	if(x==?20'b??????11???1???1?0?0) z |= 4'b0001; 
	if(x==?20'b?????????1?1??110??0) z |= 4'b0001; 
	if(x==?20'b??????1????1??110??0) z |= 4'b0001; 
	if(x==?20'b???????1??1??1?10??0) z |= 4'b0001; 
	if(x==?20'b11??1????11????????0) z |= 4'b1000; 
	if(x==?20'b1?1??1??1?1????????0) z |= 4'b1000; 
	if(x==?20'b11??1?1???1????????0) z |= 4'b1000; 
	if(x==?20'b1???1?1?11?????????0) z |= 4'b1000; 
	if(x==?20'b11????1?11?????????0) z |= 4'b1000; 
	if(x==?20'b1?1?1?1??1?????????0) z |= 4'b1000; 
	if(x==?20'b111???1??1?????????0) z |= 4'b1000; 
	if(x==?20'b???1?1?1??11???????0) z |= 4'b0100; 
	if(x==?20'b??11?1????11???????0) z |= 4'b0100; 
	if(x==?20'b?1?1??1??1?1???????0) z |= 4'b0100; 
	if(x==?20'b??11???1?11????????0) z |= 4'b0100; 
	if(x==?20'b?1?1?1?1??1????????0) z |= 4'b0100; 
	if(x==?20'b?111?1????1????????0) z |= 4'b0100; 
	if(x==?20'b??11?1?1?1?????????0) z |= 4'b0100; 
	if(x==?20'b?????1????1?111????0) z |= 4'b0010; 
	if(x==?20'b?????1??1?1?1?1????0) z |= 4'b0010; 
	if(x==?20'b????1?1??1??1?1????0) z |= 4'b0010; 
	if(x==?20'b??????1?1?1?11?????0) z |= 4'b0010; 
	if(x==?20'b????11????1?11?????0) z |= 4'b0010; 
	if(x==?20'b?????11?1???11?????0) z |= 4'b0010; 
	if(x==?20'b????11??1?1?1??????0) z |= 4'b0010; 
	if(x==?20'b??????1??1???111???0) z |= 4'b0001; 
	if(x==?20'b?????1???1?1??11???0) z |= 4'b0001; 
	if(x==?20'b?????11????1??11???0) z |= 4'b0001; 
	if(x==?20'b??????11?1????11???0) z |= 4'b0001; 
	if(x==?20'b??????1??1?1?1?1???0) z |= 4'b0001; 
	if(x==?20'b?????1?1??1??1?1???0) z |= 4'b0001; 
	if(x==?20'b??????11?1?1???1???0) z |= 4'b0001; 
	if(x==?20'b?1???1???11?????000?) z |= 4'b1000; 
	if(x==?20'b????111???1?????000?) z |= 4'b1000; 
	if(x==?20'b??1???1??11?????000?) z |= 4'b0100; 
	if(x==?20'b?????111?1??????000?) z |= 4'b0100; 
	if(x==?20'b?????11??1???1??000?) z |= 4'b0010; 
	if(x==?20'b??????1?111?????000?) z |= 4'b0010; 
	if(x==?20'b?????11???1???1?000?) z |= 4'b0001; 
	if(x==?20'b?????1???111????000?) z |= 4'b0001; 
	if(x==?20'b?????11?111??????00?) z |= 4'b1000; 
	if(x==?20'b??1??11??11??????00?) z |= 4'b1000; 
	if(x==?20'b????111??11?????0?0?) z |= 4'b1000; 
	if(x==?20'b?1???11??11?????0?0?) z |= 4'b1000; 
	if(x==?20'b?????11??111?????00?) z |= 4'b0100; 
	if(x==?20'b?1???11??11??????00?) z |= 4'b0100; 
	if(x==?20'b?????111?11?????0?0?) z |= 4'b0100; 
	if(x==?20'b??1??11??11?????0?0?) z |= 4'b0100; 
	if(x==?20'b?????11??11???1??00?) z |= 4'b0010; 
	if(x==?20'b????111??11??????00?) z |= 4'b0010; 
	if(x==?20'b?????11??11??1??0?0?) z |= 4'b0010; 
	if(x==?20'b?????11?111?????0?0?) z |= 4'b0010; 
	if(x==?20'b?????11??11??1???00?) z |= 4'b0001; 
	if(x==?20'b?????111?11??????00?) z |= 4'b0001; 
	if(x==?20'b?????11??11???1?0?0?) z |= 4'b0001; 
	if(x==?20'b?????11??111????0?0?) z |= 4'b0001; 
	if(x==?20'b?11??11?????????000?) z |= 4'b1100; 
	if(x==?20'b????11??11??????000?) z |= 4'b1010; 
	if(x==?20'b??????11??11????000?) z |= 4'b0101; 
	if(x==?20'b?????????11??11?000?) z |= 4'b0011; 
	if(x==?20'b?11??11??11???????0?) z |= 4'b1100; 
	if(x==?20'b????111?111???????0?) z |= 4'b1010; 
	if(x==?20'b?????111?111??????0?) z |= 4'b0101; 
	if(x==?20'b?????11??11??11???0?) z |= 4'b0011; 
	if(x==?20'b?1??1???1???????00?0) z |= 4'b1000; 
	if(x==?20'b?11?1???????????00?0) z |= 4'b1000; 
	if(x==?20'b??1????1???1????00?0) z |= 4'b0100; 
	if(x==?20'b?11????1????????00?0) z |= 4'b0100; 
	if(x==?20'b????????1????11?00?0) z |= 4'b0010; 
	if(x==?20'b????1???1????1??00?0) z |= 4'b0010; 
	if(x==?20'b???????????1?11?00?0) z |= 4'b0001; 
	if(x==?20'b???????1???1??1?00?0) z |= 4'b0001; 
	if(x==?20'b?1??1???1?1??????0?0) z |= 4'b1000; 
	if(x==?20'b?11?1?????1??????0?0) z |= 4'b1000; 
	if(x==?20'b??1?1???11???????0?0) z |= 4'b1000; 
	if(x==?20'b?11?????11???????0?0) z |= 4'b1000; 
	if(x==?20'b??1?1?1?1????????0?0) z |= 4'b1000; 
	if(x==?20'b?11???1?1????????0?0) z |= 4'b1000; 
	if(x==?20'b?1??1???11??????0??0) z |= 4'b1000; 
	if(x==?20'b?11?1????1??????0??0) z |= 4'b1000; 
	if(x==?20'b?1??1?1?1???????0??0) z |= 4'b1000; 
	if(x==?20'b?11?1?1?????????0??0) z |= 4'b1000; 
	if(x==?20'b?1?????1??11?????0?0) z |= 4'b0100; 
	if(x==?20'b?11???????11?????0?0) z |= 4'b0100; 
	if(x==?20'b??1????1?1?1?????0?0) z |= 4'b0100; 
	if(x==?20'b?1???1?1???1?????0?0) z |= 4'b0100; 
	if(x==?20'b?11??1?????1?????0?0) z |= 4'b0100; 
	if(x==?20'b?11????1?1???????0?0) z |= 4'b0100; 
	if(x==?20'b??1????1??11????0??0) z |= 4'b0100; 
	if(x==?20'b??1??1?1???1????0??0) z |= 4'b0100; 
	if(x==?20'b?11????1??1?????0??0) z |= 4'b0100; 
	if(x==?20'b?11??1?1????????0??0) z |= 4'b0100; 
	if(x==?20'b????1?????1??11??0?0) z |= 4'b0010; 
	if(x==?20'b??????1?1????11??0?0) z |= 4'b0010; 
	if(x==?20'b????11???????11??0?0) z |= 4'b0010; 
	if(x==?20'b????1???1?1???1??0?0) z |= 4'b0010; 
	if(x==?20'b????11??1?????1??0?0) z |= 4'b0010; 
	if(x==?20'b????1?1?1????1???0?0) z |= 4'b0010; 
	if(x==?20'b????????1?1??11?0??0) z |= 4'b0010; 
	if(x==?20'b?????1??1????11?0??0) z |= 4'b0010; 
	if(x==?20'b????1???1?1??1??0??0) z |= 4'b0010; 
	if(x==?20'b????11??1????1??0??0) z |= 4'b0010; 
	if(x==?20'b?????1?????1?11??0?0) z |= 4'b0001; 
	if(x==?20'b???????1?1???11??0?0) z |= 4'b0001; 
	if(x==?20'b??????11?????11??0?0) z |= 4'b0001; 
	if(x==?20'b?????1?1???1??1??0?0) z |= 4'b0001; 
	if(x==?20'b???????1?1?1?1???0?0) z |= 4'b0001; 
	if(x==?20'b??????11???1?1???0?0) z |= 4'b0001; 
	if(x==?20'b?????????1?1?11?0??0) z |= 4'b0001; 
	if(x==?20'b??????1????1?11?0??0) z |= 4'b0001; 
	if(x==?20'b???????1?1?1??1?0??0) z |= 4'b0001; 
	if(x==?20'b??????11???1??1?0??0) z |= 4'b0001; 
	if(x==?20'b?1??1???111????????0) z |= 4'b1000; 
	if(x==?20'b?11?1????11????????0) z |= 4'b1000; 
	if(x==?20'b?1??1?1?1?1????????0) z |= 4'b1000; 
	if(x==?20'b?11?1?1???1????????0) z |= 4'b1000; 
	if(x==?20'b??1?1?1?11?????????0) z |= 4'b1000; 
	if(x==?20'b?11???1?11?????????0) z |= 4'b1000; 
	if(x==?20'b??1????1?111???????0) z |= 4'b0100; 
	if(x==?20'b?1???1?1??11???????0) z |= 4'b0100; 
	if(x==?20'b?11??1????11???????0) z |= 4'b0100; 
	if(x==?20'b??1??1?1?1?1???????0) z |= 4'b0100; 
	if(x==?20'b?11????1?11????????0) z |= 4'b0100; 
	if(x==?20'b?11??1?1?1?????????0) z |= 4'b0100; 
	if(x==?20'b??????1?1?1??11????0) z |= 4'b0010; 
	if(x==?20'b????11????1??11????0) z |= 4'b0010; 
	if(x==?20'b?????11?1????11????0) z |= 4'b0010; 
	if(x==?20'b????11??1?1???1????0) z |= 4'b0010; 
	if(x==?20'b????1?1?1?1??1?????0) z |= 4'b0010; 
	if(x==?20'b????111?1????1?????0) z |= 4'b0010; 
	if(x==?20'b?????1???1?1?11????0) z |= 4'b0001; 
	if(x==?20'b?????11????1?11????0) z |= 4'b0001; 
	if(x==?20'b??????11?1???11????0) z |= 4'b0001; 
	if(x==?20'b?????1?1?1?1??1????0) z |= 4'b0001; 
	if(x==?20'b?????111???1??1????0) z |= 4'b0001; 
	if(x==?20'b??????11?1?1?1?????0) z |= 4'b0001; 
	if(x==?20'b1???????1?1?????0?00) z |= 4'b1000; 
	if(x==?20'b1?1???????1?????0?00) z |= 4'b1000; 
	if(x==?20'b???1?????1?1????0?00) z |= 4'b0100; 
	if(x==?20'b?1?1?????1??????0?00) z |= 4'b0100; 
	if(x==?20'b??????1?????1?1?0?00) z |= 4'b0010; 
	if(x==?20'b????1?1?????1???0?00) z |= 4'b0010; 
	if(x==?20'b?????1???????1?10?00) z |= 4'b0001; 
	if(x==?20'b?????1?1???????10?00) z |= 4'b0001; 
	if(x==?20'b1???1????1??????00?0) z |= 4'b1000; 
	if(x==?20'b11???????1??????00?0) z |= 4'b1000; 
	if(x==?20'b1???1?1?????????00?0) z |= 4'b1000; 
	if(x==?20'b11????1?????????00?0) z |= 4'b1000; 
	if(x==?20'b???1???1??1?????00?0) z |= 4'b0100; 
	if(x==?20'b??11??????1?????00?0) z |= 4'b0100; 
	if(x==?20'b???1?1?1????????00?0) z |= 4'b0100; 
	if(x==?20'b??11?1??????????00?0) z |= 4'b0100; 
	if(x==?20'b??????????1?11??00?0) z |= 4'b0010; 
	if(x==?20'b?????1??????11??00?0) z |= 4'b0010; 
	if(x==?20'b????????1?1?1???00?0) z |= 4'b0010; 
	if(x==?20'b?????1??1???1???00?0) z |= 4'b0010; 
	if(x==?20'b?????????1????1100?0) z |= 4'b0001; 
	if(x==?20'b??????1???????1100?0) z |= 4'b0001; 
	if(x==?20'b?????????1?1???100?0) z |= 4'b0001; 
	if(x==?20'b??????1????1???100?0) z |= 4'b0001; 
	if(x==?20'b1???1????11??????0?0) z |= 4'b1000; 
	if(x==?20'b11???????11??????0?0) z |= 4'b1000; 
	if(x==?20'b1???1?1???1??????0?0) z |= 4'b1000; 
	if(x==?20'b11????1???1??????0?0) z |= 4'b1000; 
	if(x==?20'b1?????1?11???????0?0) z |= 4'b1000; 
	if(x==?20'b1?1???1??1???????0?0) z |= 4'b1000; 
	if(x==?20'b1????1??1?1?????0??0) z |= 4'b1000; 
	if(x==?20'b1?1??1????1?????0??0) z |= 4'b1000; 
	if(x==?20'b1???1?1??1??????0??0) z |= 4'b1000; 
	if(x==?20'b11????1??1??????0??0) z |= 4'b1000; 
	if(x==?20'b???1?1????11?????0?0) z |= 4'b0100; 
	if(x==?20'b???1???1?11??????0?0) z |= 4'b0100; 
	if(x==?20'b??11?????11??????0?0) z |= 4'b0100; 
	if(x==?20'b?1?1?1????1??????0?0) z |= 4'b0100; 
	if(x==?20'b???1?1?1?1???????0?0) z |= 4'b0100; 
	if(x==?20'b??11?1???1???????0?0) z |= 4'b0100; 
	if(x==?20'b???1??1??1?1????0??0) z |= 4'b0100; 
	if(x==?20'b???1?1?1??1?????0??0) z |= 4'b0100; 
	if(x==?20'b??11?1????1?????0??0) z |= 4'b0100; 
	if(x==?20'b?1?1??1??1??????0??0) z |= 4'b0100; 
	if(x==?20'b?????1????1?1?1??0?0) z |= 4'b0010; 
	if(x==?20'b??????1???1?11???0?0) z |= 4'b0010; 
	if(x==?20'b?????11?????11???0?0) z |= 4'b0010; 
	if(x==?20'b??????1?1?1?1????0?0) z |= 4'b0010; 
	if(x==?20'b????11????1?1????0?0) z |= 4'b0010; 
	if(x==?20'b?????11?1???1????0?0) z |= 4'b0010; 
	if(x==?20'b??????1??1??1?1?0??0) z |= 4'b0010; 
	if(x==?20'b?????1????1?11??0??0) z |= 4'b0010; 
	if(x==?20'b?????1??1?1?1???0??0) z |= 4'b0010; 
	if(x==?20'b????1?1??1??1???0??0) z |= 4'b0010; 
	if(x==?20'b?????1???1????11?0?0) z |= 4'b0001; 
	if(x==?20'b?????11???????11?0?0) z |= 4'b0001; 
	if(x==?20'b??????1??1???1?1?0?0) z |= 4'b0001; 
	if(x==?20'b?????1???1?1???1?0?0) z |= 4'b0001; 
	if(x==?20'b?????11????1???1?0?0) z |= 4'b0001; 
	if(x==?20'b??????11?1?????1?0?0) z |= 4'b0001; 
	if(x==?20'b??????1??1????110??0) z |= 4'b0001; 
	if(x==?20'b?????1????1??1?10??0) z |= 4'b0001; 
	if(x==?20'b??????1??1?1???10??0) z |= 4'b0001; 
	if(x==?20'b?????1?1??1????10??0) z |= 4'b0001; 
	if(x==?20'b1???1?1??11????????0) z |= 4'b1000; 
	if(x==?20'b11????1??11????????0) z |= 4'b1000; 
	if(x==?20'b???1?1?1?11????????0) z |= 4'b0100; 
	if(x==?20'b??11?1???11????????0) z |= 4'b0100; 
	if(x==?20'b?????11???1?11?????0) z |= 4'b0010; 
	if(x==?20'b?????11?1?1?1??????0) z |= 4'b0010; 
	if(x==?20'b?????11??1????11???0) z |= 4'b0001; 
	if(x==?20'b?????11??1?1???1???0) z |= 4'b0001; 
	if(x==?20'b?1??11???1???????00?) z |= 4'b1000; 
	if(x==?20'b?1??111??????????00?) z |= 4'b1000; 
	if(x==?20'b??1???11??1??????00?) z |= 4'b0100; 
	if(x==?20'b??1??111?????????00?) z |= 4'b0100; 
	if(x==?20'b????????111??1???00?) z |= 4'b0010; 
	if(x==?20'b?????1??11???1???00?) z |= 4'b0010; 
	if(x==?20'b?????????111??1??00?) z |= 4'b0001; 
	if(x==?20'b??????1???11??1??00?) z |= 4'b0001; 
	if(x==?20'b?1???11???1?????000?) z |= 4'b1100; 
	if(x==?20'b??1??11??1??????000?) z |= 4'b1100; 
	if(x==?20'b????11???11?????000?) z |= 4'b1010; 
	if(x==?20'b?????11?11??????000?) z |= 4'b1010; 
	if(x==?20'b?????11???11????000?) z |= 4'b0101; 
	if(x==?20'b??????11?11?????000?) z |= 4'b0101; 
	if(x==?20'b?????1???11???1?000?) z |= 4'b0011; 
	if(x==?20'b??????1??11??1??000?) z |= 4'b0011; 
	if(x==?20'b?1??111??1????????0?) z |= 4'b1000; 
	if(x==?20'b??1??111??1???????0?) z |= 4'b0100; 
	if(x==?20'b?????1??111??1????0?) z |= 4'b0010; 
	if(x==?20'b??????1??111??1???0?) z |= 4'b0001; 
	if(x==?20'b??1?????1?1?????0?00) z |= 4'b1000; 
	if(x==?20'b?1???????1?1????0?00) z |= 4'b0100; 
	if(x==?20'b????1?1???????1?0?00) z |= 4'b0010; 
	if(x==?20'b?????1?1?????1??0?00) z |= 4'b0001; 
	if(x==?20'b?1??1?????1?????00?0) z |= 4'b1000; 
	if(x==?20'b????1???11??????00?0) z |= 4'b1000; 
	if(x==?20'b?1??????11??????00?0) z |= 4'b1000; 
	if(x==?20'b??1?1????1??????00?0) z |= 4'b1000; 
	if(x==?20'b?11??????1??????00?0) z |= 4'b1000; 
	if(x==?20'b????1?1?1???????00?0) z |= 4'b1000; 
	if(x==?20'b?1????1?1???????00?0) z |= 4'b1000; 
	if(x==?20'b??1?1?1?????????00?0) z |= 4'b1000; 
	if(x==?20'b?11???1?????????00?0) z |= 4'b1000; 
	if(x==?20'b???????1??11????00?0) z |= 4'b0100; 
	if(x==?20'b??1???????11????00?0) z |= 4'b0100; 
	if(x==?20'b?????1?1???1????00?0) z |= 4'b0100; 
	if(x==?20'b??1??1?????1????00?0) z |= 4'b0100; 
	if(x==?20'b?1?????1??1?????00?0) z |= 4'b0100; 
	if(x==?20'b?11???????1?????00?0) z |= 4'b0100; 
	if(x==?20'b??1????1?1??????00?0) z |= 4'b0100; 
	if(x==?20'b?1???1?1????????00?0) z |= 4'b0100; 
	if(x==?20'b?11??1??????????00?0) z |= 4'b0100; 
	if(x==?20'b??????????1??11?00?0) z |= 4'b0010; 
	if(x==?20'b?????1???????11?00?0) z |= 4'b0010; 
	if(x==?20'b????????1?1???1?00?0) z |= 4'b0010; 
	if(x==?20'b?????1??1?????1?00?0) z |= 4'b0010; 
	if(x==?20'b????1?????1??1??00?0) z |= 4'b0010; 
	if(x==?20'b??????1?1????1??00?0) z |= 4'b0010; 
	if(x==?20'b????11???????1??00?0) z |= 4'b0010; 
	if(x==?20'b????1???1?1?????00?0) z |= 4'b0010; 
	if(x==?20'b????11??1???????00?0) z |= 4'b0010; 
	if(x==?20'b?????????1???11?00?0) z |= 4'b0001; 
	if(x==?20'b??????1??????11?00?0) z |= 4'b0001; 
	if(x==?20'b?????1?????1??1?00?0) z |= 4'b0001; 
	if(x==?20'b???????1?1????1?00?0) z |= 4'b0001; 
	if(x==?20'b??????11??????1?00?0) z |= 4'b0001; 
	if(x==?20'b?????????1?1?1??00?0) z |= 4'b0001; 
	if(x==?20'b??????1????1?1??00?0) z |= 4'b0001; 
	if(x==?20'b???????1?1?1????00?0) z |= 4'b0001; 
	if(x==?20'b??????11???1????00?0) z |= 4'b0001; 
	if(x==?20'b????1???111??????0?0) z |= 4'b1000; 
	if(x==?20'b?1??????111??????0?0) z |= 4'b1000; 
	if(x==?20'b??1?1????11??????0?0) z |= 4'b1000; 
	if(x==?20'b?1????1?1?1??????0?0) z |= 4'b1000; 
	if(x==?20'b??1?1?1???1??????0?0) z |= 4'b1000; 
	if(x==?20'b?11???1???1??????0?0) z |= 4'b1000; 
	if(x==?20'b??1???1?11???????0?0) z |= 4'b1000; 
	if(x==?20'b?1??1????11?????0??0) z |= 4'b1000; 
	if(x==?20'b??1??1??1?1?????0??0) z |= 4'b1000; 
	if(x==?20'b?1??1?1???1?????0??0) z |= 4'b1000; 
	if(x==?20'b????1?1?11??????0??0) z |= 4'b1000; 
	if(x==?20'b?1????1?11??????0??0) z |= 4'b1000; 
	if(x==?20'b??1?1?1??1??????0??0) z |= 4'b1000; 
	if(x==?20'b?11???1??1??????0??0) z |= 4'b1000; 
	if(x==?20'b???????1?111?????0?0) z |= 4'b0100; 
	if(x==?20'b??1??????111?????0?0) z |= 4'b0100; 
	if(x==?20'b?1???1????11?????0?0) z |= 4'b0100; 
	if(x==?20'b??1??1???1?1?????0?0) z |= 4'b0100; 
	if(x==?20'b?1?????1?11??????0?0) z |= 4'b0100; 
	if(x==?20'b?1???1?1?1???????0?0) z |= 4'b0100; 
	if(x==?20'b?11??1???1???????0?0) z |= 4'b0100; 
	if(x==?20'b?????1?1??11????0??0) z |= 4'b0100; 
	if(x==?20'b??1??1????11????0??0) z |= 4'b0100; 
	if(x==?20'b?1????1??1?1????0??0) z |= 4'b0100; 
	if(x==?20'b??1????1?11?????0??0) z |= 4'b0100; 
	if(x==?20'b?1???1?1??1?????0??0) z |= 4'b0100; 
	if(x==?20'b?11??1????1?????0??0) z |= 4'b0100; 
	if(x==?20'b??1??1?1?1??????0??0) z |= 4'b0100; 
	if(x==?20'b??????1???1??11??0?0) z |= 4'b0010; 
	if(x==?20'b??????1?1?1???1??0?0) z |= 4'b0010; 
	if(x==?20'b????11????1???1??0?0) z |= 4'b0010; 
	if(x==?20'b?????11?1?????1??0?0) z |= 4'b0010; 
	if(x==?20'b????1?1???1??1???0?0) z |= 4'b0010; 
	if(x==?20'b????111??????1???0?0) z |= 4'b0010; 
	if(x==?20'b????111?1????????0?0) z |= 4'b0010; 
	if(x==?20'b?????1????1??11?0??0) z |= 4'b0010; 
	if(x==?20'b?????1??1?1???1?0??0) z |= 4'b0010; 
	if(x==?20'b????1?1??1????1?0??0) z |= 4'b0010; 
	if(x==?20'b??????1?1?1??1??0??0) z |= 4'b0010; 
	if(x==?20'b????11????1??1??0??0) z |= 4'b0010; 
	if(x==?20'b?????11?1????1??0??0) z |= 4'b0010; 
	if(x==?20'b????11??1?1?????0??0) z |= 4'b0010; 
	if(x==?20'b?????1???1???11??0?0) z |= 4'b0001; 
	if(x==?20'b?????1?1?1????1??0?0) z |= 4'b0001; 
	if(x==?20'b?????111??????1??0?0) z |= 4'b0001; 
	if(x==?20'b?????1???1?1?1???0?0) z |= 4'b0001; 
	if(x==?20'b?????11????1?1???0?0) z |= 4'b0001; 
	if(x==?20'b??????11?1???1???0?0) z |= 4'b0001; 
	if(x==?20'b?????111???1?????0?0) z |= 4'b0001; 
	if(x==?20'b??????1??1???11?0??0) z |= 4'b0001; 
	if(x==?20'b?????1???1?1??1?0??0) z |= 4'b0001; 
	if(x==?20'b?????11????1??1?0??0) z |= 4'b0001; 
	if(x==?20'b??????11?1????1?0??0) z |= 4'b0001; 
	if(x==?20'b??????1??1?1?1??0??0) z |= 4'b0001; 
	if(x==?20'b?????1?1??1??1??0??0) z |= 4'b0001; 
	if(x==?20'b??????11?1?1????0??0) z |= 4'b0001; 
	if(x==?20'b????1?1?111????????0) z |= 4'b1000; 
	if(x==?20'b?1????1?111????????0) z |= 4'b1000; 
	if(x==?20'b??1?1?1??11????????0) z |= 4'b1000; 
	if(x==?20'b?11???1??11????????0) z |= 4'b1000; 
	if(x==?20'b?????1?1?111???????0) z |= 4'b0100; 
	if(x==?20'b??1??1???111???????0) z |= 4'b0100; 
	if(x==?20'b?1???1?1?11????????0) z |= 4'b0100; 
	if(x==?20'b?11??1???11????????0) z |= 4'b0100; 
	if(x==?20'b?????11???1??11????0) z |= 4'b0010; 
	if(x==?20'b?????11?1?1???1????0) z |= 4'b0010; 
	if(x==?20'b????111???1??1?????0) z |= 4'b0010; 
	if(x==?20'b????111?1?1????????0) z |= 4'b0010; 
	if(x==?20'b?????11??1???11????0) z |= 4'b0001; 
	if(x==?20'b?????111?1????1????0) z |= 4'b0001; 
	if(x==?20'b?????11??1?1?1?????0) z |= 4'b0001; 
	if(x==?20'b?????111?1?1???????0) z |= 4'b0001; 
	if(x==?20'b1?????1??1??????00?0) z |= 4'b1000; 
	if(x==?20'b???1?1????1?????00?0) z |= 4'b0100; 
	if(x==?20'b?????1????1?1???00?0) z |= 4'b0010; 
	if(x==?20'b??????1??1?????100?0) z |= 4'b0001; 
	if(x==?20'b1?????1??11??????0?0) z |= 4'b1000; 
	if(x==?20'b???1?1???11??????0?0) z |= 4'b0100; 
	if(x==?20'b?????11???1?1????0?0) z |= 4'b0010; 
	if(x==?20'b?????11??1?????1?0?0) z |= 4'b0001; 
	if(x==?20'b1???1???1?????????00) z |= 4'b1000; 
	if(x==?20'b11??????1?????????00) z |= 4'b1000; 
	if(x==?20'b1?1?1?????????????00) z |= 4'b1000; 
	if(x==?20'b111???????????????00) z |= 4'b1000; 
	if(x==?20'b???1???1???1??????00) z |= 4'b0100; 
	if(x==?20'b??11???????1??????00) z |= 4'b0100; 
	if(x==?20'b?1?1???1??????????00) z |= 4'b0100; 
	if(x==?20'b?111??????????????00) z |= 4'b0100; 
	if(x==?20'b????????????111???00) z |= 4'b0010; 
	if(x==?20'b????????1???1?1???00) z |= 4'b0010; 
	if(x==?20'b????1???????11????00) z |= 4'b0010; 
	if(x==?20'b????1???1???1?????00) z |= 4'b0010; 
	if(x==?20'b?????????????111??00) z |= 4'b0001; 
	if(x==?20'b???????1??????11??00) z |= 4'b0001; 
	if(x==?20'b???????????1?1?1??00) z |= 4'b0001; 
	if(x==?20'b???????1???1???1??00) z |= 4'b0001; 
	if(x==?20'b1???11??1??????????0) z |= 4'b1000; 
	if(x==?20'b11???1??1??????????0) z |= 4'b1000; 
	if(x==?20'b1?1?11?????????????0) z |= 4'b1000; 
	if(x==?20'b111??1?????????????0) z |= 4'b1000; 
	if(x==?20'b???1??11???1???????0) z |= 4'b0100; 
	if(x==?20'b??11??1????1???????0) z |= 4'b0100; 
	if(x==?20'b?1?1??11???????????0) z |= 4'b0100; 
	if(x==?20'b?111??1????????????0) z |= 4'b0100; 
	if(x==?20'b?????????1??111????0) z |= 4'b0010; 
	if(x==?20'b????????11??1?1????0) z |= 4'b0010; 
	if(x==?20'b????1????1??11?????0) z |= 4'b0010; 
	if(x==?20'b????1???11??1??????0) z |= 4'b0010; 
	if(x==?20'b??????????1??111???0) z |= 4'b0001; 
	if(x==?20'b???????1??1???11???0) z |= 4'b0001; 
	if(x==?20'b??????????11?1?1???0) z |= 4'b0001; 
	if(x==?20'b???????1??11???1???0) z |= 4'b0001; 
	if(x==?20'b????111??1???????00?) z |= 4'b1000; 
	if(x==?20'b?1???11??1???????00?) z |= 4'b1000; 
	if(x==?20'b?????111??1??????00?) z |= 4'b0100; 
	if(x==?20'b??1??11???1??????00?) z |= 4'b0100; 
	if(x==?20'b?????1???11??1???00?) z |= 4'b0010; 
	if(x==?20'b?????1??111??????00?) z |= 4'b0010; 
	if(x==?20'b??????1??11???1??00?) z |= 4'b0001; 
	if(x==?20'b??????1??111?????00?) z |= 4'b0001; 
	if(x==?20'b????1????11?????00?0) z |= 4'b1000; 
	if(x==?20'b?1???????11?????00?0) z |= 4'b1000; 
	if(x==?20'b????1?1???1?????00?0) z |= 4'b1000; 
	if(x==?20'b?1????1???1?????00?0) z |= 4'b1000; 
	if(x==?20'b??????1?11??????00?0) z |= 4'b1000; 
	if(x==?20'b??1???1??1??????00?0) z |= 4'b1000; 
	if(x==?20'b?????1????11????00?0) z |= 4'b0100; 
	if(x==?20'b???????1?11?????00?0) z |= 4'b0100; 
	if(x==?20'b??1??????11?????00?0) z |= 4'b0100; 
	if(x==?20'b?1???1????1?????00?0) z |= 4'b0100; 
	if(x==?20'b?????1?1?1??????00?0) z |= 4'b0100; 
	if(x==?20'b??1??1???1??????00?0) z |= 4'b0100; 
	if(x==?20'b?????1????1???1?00?0) z |= 4'b0010; 
	if(x==?20'b??????1???1??1??00?0) z |= 4'b0010; 
	if(x==?20'b?????11??????1??00?0) z |= 4'b0010; 
	if(x==?20'b??????1?1?1?????00?0) z |= 4'b0010; 
	if(x==?20'b????11????1?????00?0) z |= 4'b0010; 
	if(x==?20'b?????11?1???????00?0) z |= 4'b0010; 
	if(x==?20'b?????1???1????1?00?0) z |= 4'b0001; 
	if(x==?20'b?????11???????1?00?0) z |= 4'b0001; 
	if(x==?20'b??????1??1???1??00?0) z |= 4'b0001; 
	if(x==?20'b?????1???1?1????00?0) z |= 4'b0001; 
	if(x==?20'b?????11????1????00?0) z |= 4'b0001; 
	if(x==?20'b??????11?1??????00?0) z |= 4'b0001; 
	if(x==?20'b??????1?111??????0?0) z |= 4'b1000; 
	if(x==?20'b??1???1??11??????0?0) z |= 4'b1000; 
	if(x==?20'b????1?1??11?????0??0) z |= 4'b1000; 
	if(x==?20'b?1????1??11?????0??0) z |= 4'b1000; 
	if(x==?20'b?????1???111?????0?0) z |= 4'b0100; 
	if(x==?20'b?1???1???11??????0?0) z |= 4'b0100; 
	if(x==?20'b?????1?1?11?????0??0) z |= 4'b0100; 
	if(x==?20'b??1??1???11?????0??0) z |= 4'b0100; 
	if(x==?20'b?????11???1???1??0?0) z |= 4'b0010; 
	if(x==?20'b????111???1??????0?0) z |= 4'b0010; 
	if(x==?20'b?????11???1??1??0??0) z |= 4'b0010; 
	if(x==?20'b?????11?1?1?????0??0) z |= 4'b0010; 
	if(x==?20'b?????11??1???1???0?0) z |= 4'b0001; 
	if(x==?20'b?????111?1???????0?0) z |= 4'b0001; 
	if(x==?20'b?????11??1????1?0??0) z |= 4'b0001; 
	if(x==?20'b?????11??1?1????0??0) z |= 4'b0001; 
	if(x==?20'b??1?1???1?????????00) z |= 4'b1000; 
	if(x==?20'b?11?????1?????????00) z |= 4'b1000; 
	if(x==?20'b?1?????1???1??????00) z |= 4'b0100; 
	if(x==?20'b?11????????1??????00) z |= 4'b0100; 
	if(x==?20'b????1????????11???00) z |= 4'b0010; 
	if(x==?20'b????1???1?????1???00) z |= 4'b0010; 
	if(x==?20'b???????1?????11???00) z |= 4'b0001; 
	if(x==?20'b???????1???1?1????00) z |= 4'b0001; 
	if(x==?20'b??1?11??1??????????0) z |= 4'b1000; 
	if(x==?20'b?11??1??1??????????0) z |= 4'b1000; 
	if(x==?20'b?1????11???1???????0) z |= 4'b0100; 
	if(x==?20'b?11???1????1???????0) z |= 4'b0100; 
	if(x==?20'b????1????1???11????0) z |= 4'b0010; 
	if(x==?20'b????1???11????1????0) z |= 4'b0010; 
	if(x==?20'b???????1??1??11????0) z |= 4'b0001; 
	if(x==?20'b???????1??11?1?????0) z |= 4'b0001; 
	if(x==?20'b?11??????11??????0?0) z |= 4'b1100; 
	if(x==?20'b????1?1?1?1??????0?0) z |= 4'b1010; 
	if(x==?20'b?????1?1?1?1?????0?0) z |= 4'b0101; 
	if(x==?20'b?????11??????11??0?0) z |= 4'b0011; 
	if(x==?20'b1???????1????????000) z |= 4'b1000; 
	if(x==?20'b1?1??????????????000) z |= 4'b1000; 
	if(x==?20'b1???1???????????0?00) z |= 4'b1000; 
	if(x==?20'b11??????????????0?00) z |= 4'b1000; 
	if(x==?20'b???1???????1?????000) z |= 4'b0100; 
	if(x==?20'b?1?1?????????????000) z |= 4'b0100; 
	if(x==?20'b???1???1????????0?00) z |= 4'b0100; 
	if(x==?20'b??11????????????0?00) z |= 4'b0100; 
	if(x==?20'b????????????1?1??000) z |= 4'b0010; 
	if(x==?20'b????1???????1????000) z |= 4'b0010; 
	if(x==?20'b????????????11??0?00) z |= 4'b0010; 
	if(x==?20'b????????1???1???0?00) z |= 4'b0010; 
	if(x==?20'b?????????????1?1?000) z |= 4'b0001; 
	if(x==?20'b???????1???????1?000) z |= 4'b0001; 
	if(x==?20'b??????????????110?00) z |= 4'b0001; 
	if(x==?20'b???????????1???10?00) z |= 4'b0001; 
	if(x==?20'b1???1?????1???????00) z |= 4'b1000; 
	if(x==?20'b11????????1???????00) z |= 4'b1000; 
	if(x==?20'b1???????11????????00) z |= 4'b1000; 
	if(x==?20'b1?1??????1????????00) z |= 4'b1000; 
	if(x==?20'b1?????1?1?????????00) z |= 4'b1000; 
	if(x==?20'b1?1???1???????????00) z |= 4'b1000; 
	if(x==?20'b???1??????11??????00) z |= 4'b0100; 
	if(x==?20'b???1?1?????1??????00) z |= 4'b0100; 
	if(x==?20'b?1?1??????1???????00) z |= 4'b0100; 
	if(x==?20'b???1???1?1????????00) z |= 4'b0100; 
	if(x==?20'b??11?????1????????00) z |= 4'b0100; 
	if(x==?20'b?1?1?1????????????00) z |= 4'b0100; 
	if(x==?20'b??????????1?1?1???00) z |= 4'b0010; 
	if(x==?20'b?????1??????1?1???00) z |= 4'b0010; 
	if(x==?20'b??????1?????11????00) z |= 4'b0010; 
	if(x==?20'b????1?????1?1?????00) z |= 4'b0010; 
	if(x==?20'b??????1?1???1?????00) z |= 4'b0010; 
	if(x==?20'b????11??????1?????00) z |= 4'b0010; 
	if(x==?20'b?????1????????11??00) z |= 4'b0001; 
	if(x==?20'b?????????1???1?1??00) z |= 4'b0001; 
	if(x==?20'b??????1??????1?1??00) z |= 4'b0001; 
	if(x==?20'b?????1?????1???1??00) z |= 4'b0001; 
	if(x==?20'b???????1?1?????1??00) z |= 4'b0001; 
	if(x==?20'b??????11???????1??00) z |= 4'b0001; 
	if(x==?20'b1????1??1????????0?0) z |= 4'b1000; 
	if(x==?20'b1?1??1???????????0?0) z |= 4'b1000; 
	if(x==?20'b1???11??????????0??0) z |= 4'b1000; 
	if(x==?20'b11???1??????????0??0) z |= 4'b1000; 
	if(x==?20'b???1??1????1?????0?0) z |= 4'b0100; 
	if(x==?20'b?1?1??1??????????0?0) z |= 4'b0100; 
	if(x==?20'b???1??11????????0??0) z |= 4'b0100; 
	if(x==?20'b??11??1?????????0??0) z |= 4'b0100; 
	if(x==?20'b?????????1??1?1??0?0) z |= 4'b0010; 
	if(x==?20'b????1????1??1????0?0) z |= 4'b0010; 
	if(x==?20'b?????????1??11??0??0) z |= 4'b0010; 
	if(x==?20'b????????11??1???0??0) z |= 4'b0010; 
	if(x==?20'b??????????1??1?1?0?0) z |= 4'b0001; 
	if(x==?20'b???????1??1????1?0?0) z |= 4'b0001; 
	if(x==?20'b??????????1???110??0) z |= 4'b0001; 
	if(x==?20'b??????????11???10??0) z |= 4'b0001; 
	if(x==?20'b1???11????1????????0) z |= 4'b1000; 
	if(x==?20'b11???1????1????????0) z |= 4'b1000; 
	if(x==?20'b1????1??11?????????0) z |= 4'b1000; 
	if(x==?20'b1?1??1???1?????????0) z |= 4'b1000; 
	if(x==?20'b1????11?1??????????0) z |= 4'b1000; 
	if(x==?20'b1?1??11????????????0) z |= 4'b1000; 
	if(x==?20'b???1??1???11???????0) z |= 4'b0100; 
	if(x==?20'b???1?11????1???????0) z |= 4'b0100; 
	if(x==?20'b?1?1??1???1????????0) z |= 4'b0100; 
	if(x==?20'b???1??11?1?????????0) z |= 4'b0100; 
	if(x==?20'b??11??1??1?????????0) z |= 4'b0100; 
	if(x==?20'b?1?1?11????????????0) z |= 4'b0100; 
	if(x==?20'b?????????11?1?1????0) z |= 4'b0010; 
	if(x==?20'b?????1???1??1?1????0) z |= 4'b0010; 
	if(x==?20'b??????1??1??11?????0) z |= 4'b0010; 
	if(x==?20'b????1????11?1??????0) z |= 4'b0010; 
	if(x==?20'b??????1?11??1??????0) z |= 4'b0010; 
	if(x==?20'b????11???1??1??????0) z |= 4'b0010; 
	if(x==?20'b?????1????1???11???0) z |= 4'b0001; 
	if(x==?20'b?????????11??1?1???0) z |= 4'b0001; 
	if(x==?20'b??????1???1??1?1???0) z |= 4'b0001; 
	if(x==?20'b?????1????11???1???0) z |= 4'b0001; 
	if(x==?20'b???????1?11????1???0) z |= 4'b0001; 
	if(x==?20'b??????11??1????1???0) z |= 4'b0001; 
	if(x==?20'b??????1??11?????00?0) z |= 4'b1000; 
	if(x==?20'b?????1???11?????00?0) z |= 4'b0100; 
	if(x==?20'b?????11???1?????00?0) z |= 4'b0010; 
	if(x==?20'b?????11??1??????00?0) z |= 4'b0001; 
	if(x==?20'b??1?????1????????000) z |= 4'b1000; 
	if(x==?20'b?1??????1???????0?00) z |= 4'b1000; 
	if(x==?20'b??1?1???????????0?00) z |= 4'b1000; 
	if(x==?20'b?1?????????1?????000) z |= 4'b0100; 
	if(x==?20'b??1????????1????0?00) z |= 4'b0100; 
	if(x==?20'b?1?????1????????0?00) z |= 4'b0100; 
	if(x==?20'b????1?????????1??000) z |= 4'b0010; 
	if(x==?20'b????????1?????1?0?00) z |= 4'b0010; 
	if(x==?20'b????1????????1??0?00) z |= 4'b0010; 
	if(x==?20'b???????1?????1???000) z |= 4'b0001; 
	if(x==?20'b???????1??????1?0?00) z |= 4'b0001; 
	if(x==?20'b???????????1?1??0?00) z |= 4'b0001; 
	if(x==?20'b????1???1?1???????00) z |= 4'b1000; 
	if(x==?20'b?1??????1?1???????00) z |= 4'b1000; 
	if(x==?20'b??1?1?????1???????00) z |= 4'b1000; 
	if(x==?20'b?11???????1???????00) z |= 4'b1000; 
	if(x==?20'b??1?????11????????00) z |= 4'b1000; 
	if(x==?20'b??1???1?1?????????00) z |= 4'b1000; 
	if(x==?20'b?1????????11??????00) z |= 4'b0100; 
	if(x==?20'b???????1?1?1??????00) z |= 4'b0100; 
	if(x==?20'b??1??????1?1??????00) z |= 4'b0100; 
	if(x==?20'b?1???1?????1??????00) z |= 4'b0100; 
	if(x==?20'b?1?????1?1????????00) z |= 4'b0100; 
	if(x==?20'b?11??????1????????00) z |= 4'b0100; 
	if(x==?20'b??????1??????11???00) z |= 4'b0010; 
	if(x==?20'b????1?????1???1???00) z |= 4'b0010; 
	if(x==?20'b??????1?1?????1???00) z |= 4'b0010; 
	if(x==?20'b????11????????1???00) z |= 4'b0010; 
	if(x==?20'b????1?1??????1????00) z |= 4'b0010; 
	if(x==?20'b????1?1?1?????????00) z |= 4'b0010; 
	if(x==?20'b?????1???????11???00) z |= 4'b0001; 
	if(x==?20'b?????1?1??????1???00) z |= 4'b0001; 
	if(x==?20'b?????1?????1?1????00) z |= 4'b0001; 
	if(x==?20'b???????1?1???1????00) z |= 4'b0001; 
	if(x==?20'b??????11?????1????00) z |= 4'b0001; 
	if(x==?20'b?????1?1???1??????00) z |= 4'b0001; 
	if(x==?20'b?1??1????1???????0?0) z |= 4'b1000; 
	if(x==?20'b??1??1??1????????0?0) z |= 4'b1000; 
	if(x==?20'b?1??1?1??????????0?0) z |= 4'b1000; 
	if(x==?20'b????11??1???????0??0) z |= 4'b1000; 
	if(x==?20'b?1???1??1???????0??0) z |= 4'b1000; 
	if(x==?20'b??1?11??????????0??0) z |= 4'b1000; 
	if(x==?20'b?11??1??????????0??0) z |= 4'b1000; 
	if(x==?20'b?1????1????1?????0?0) z |= 4'b0100; 
	if(x==?20'b??1????1??1??????0?0) z |= 4'b0100; 
	if(x==?20'b??1??1?1?????????0?0) z |= 4'b0100; 
	if(x==?20'b??????11???1????0??0) z |= 4'b0100; 
	if(x==?20'b??1???1????1????0??0) z |= 4'b0100; 
	if(x==?20'b?1????11????????0??0) z |= 4'b0100; 
	if(x==?20'b?11???1?????????0??0) z |= 4'b0100; 
	if(x==?20'b????1????1????1??0?0) z |= 4'b0010; 
	if(x==?20'b????????1?1??1???0?0) z |= 4'b0010; 
	if(x==?20'b?????1??1????1???0?0) z |= 4'b0010; 
	if(x==?20'b?????????1???11?0??0) z |= 4'b0010; 
	if(x==?20'b????????11????1?0??0) z |= 4'b0010; 
	if(x==?20'b????1????1???1??0??0) z |= 4'b0010; 
	if(x==?20'b????1???11??????0??0) z |= 4'b0010; 
	if(x==?20'b?????????1?1??1??0?0) z |= 4'b0001; 
	if(x==?20'b??????1????1??1??0?0) z |= 4'b0001; 
	if(x==?20'b???????1??1??1???0?0) z |= 4'b0001; 
	if(x==?20'b??????????1??11?0??0) z |= 4'b0001; 
	if(x==?20'b???????1??1???1?0??0) z |= 4'b0001; 
	if(x==?20'b??????????11?1??0??0) z |= 4'b0001; 
	if(x==?20'b???????1??11????0??0) z |= 4'b0001; 
	if(x==?20'b????11??1?1????????0) z |= 4'b1000; 
	if(x==?20'b?1???1??1?1????????0) z |= 4'b1000; 
	if(x==?20'b??1?11????1????????0) z |= 4'b1000; 
	if(x==?20'b?11??1????1????????0) z |= 4'b1000; 
	if(x==?20'b??1??1??11?????????0) z |= 4'b1000; 
	if(x==?20'b?1??1?1??1?????????0) z |= 4'b1000; 
	if(x==?20'b??1??11?1??????????0) z |= 4'b1000; 
	if(x==?20'b?1????1???11???????0) z |= 4'b0100; 
	if(x==?20'b??????11?1?1???????0) z |= 4'b0100; 
	if(x==?20'b??1???1??1?1???????0) z |= 4'b0100; 
	if(x==?20'b?1???11????1???????0) z |= 4'b0100; 
	if(x==?20'b??1??1?1??1????????0) z |= 4'b0100; 
	if(x==?20'b?1????11?1?????????0) z |= 4'b0100; 
	if(x==?20'b?11???1??1?????????0) z |= 4'b0100; 
	if(x==?20'b??????1??1???11????0) z |= 4'b0010; 
	if(x==?20'b????1????11???1????0) z |= 4'b0010; 
	if(x==?20'b??????1?11????1????0) z |= 4'b0010; 
	if(x==?20'b????11???1????1????0) z |= 4'b0010; 
	if(x==?20'b?????1??1?1??1?????0) z |= 4'b0010; 
	if(x==?20'b????1?1??1???1?????0) z |= 4'b0010; 
	if(x==?20'b????1?1?11?????????0) z |= 4'b0010; 
	if(x==?20'b?????1????1??11????0) z |= 4'b0001; 
	if(x==?20'b??????1??1?1??1????0) z |= 4'b0001; 
	if(x==?20'b?????1?1??1???1????0) z |= 4'b0001; 
	if(x==?20'b?????1????11?1?????0) z |= 4'b0001; 
	if(x==?20'b???????1?11??1?????0) z |= 4'b0001; 
	if(x==?20'b??????11??1??1?????0) z |= 4'b0001; 
	if(x==?20'b?????1?1??11???????0) z |= 4'b0001; 
	if(x==?20'b1???????????????0000) z |= 4'b1000; 
	if(x==?20'b???1????????????0000) z |= 4'b0100; 
	if(x==?20'b????????????1???0000) z |= 4'b0010; 
	if(x==?20'b???????????????10000) z |= 4'b0001; 
	if(x==?20'b1?????????1??????000) z |= 4'b1000; 
	if(x==?20'b1????????1??????0?00) z |= 4'b1000; 
	if(x==?20'b1?????1?????????0?00) z |= 4'b1000; 
	if(x==?20'b???1?????1???????000) z |= 4'b0100; 
	if(x==?20'b???1??????1?????0?00) z |= 4'b0100; 
	if(x==?20'b???1?1??????????0?00) z |= 4'b0100; 
	if(x==?20'b??????1?????1????000) z |= 4'b0010; 
	if(x==?20'b??????????1?1???0?00) z |= 4'b0010; 
	if(x==?20'b?????1??????1???0?00) z |= 4'b0010; 
	if(x==?20'b?????1?????????1?000) z |= 4'b0001; 
	if(x==?20'b?????????1?????10?00) z |= 4'b0001; 
	if(x==?20'b??????1????????10?00) z |= 4'b0001; 
	if(x==?20'b1????????11???????00) z |= 4'b1000; 
	if(x==?20'b1?????1???1???????00) z |= 4'b1000; 
	if(x==?20'b1????1??????????00?0) z |= 4'b1000; 
	if(x==?20'b???1?????11???????00) z |= 4'b0100; 
	if(x==?20'b???1?1???1????????00) z |= 4'b0100; 
	if(x==?20'b???1??1?????????00?0) z |= 4'b0100; 
	if(x==?20'b??????1???1?1?????00) z |= 4'b0010; 
	if(x==?20'b?????11?????1?????00) z |= 4'b0010; 
	if(x==?20'b?????????1??1???00?0) z |= 4'b0010; 
	if(x==?20'b?????1???1?????1??00) z |= 4'b0001; 
	if(x==?20'b?????11????????1??00) z |= 4'b0001; 
	if(x==?20'b??????????1????100?0) z |= 4'b0001; 
	if(x==?20'b1????1????1??????0?0) z |= 4'b1000; 
	if(x==?20'b1????1???1??????0??0) z |= 4'b1000; 
	if(x==?20'b1????11?????????0??0) z |= 4'b1000; 
	if(x==?20'b???1??1??1???????0?0) z |= 4'b0100; 
	if(x==?20'b???1??1???1?????0??0) z |= 4'b0100; 
	if(x==?20'b???1?11?????????0??0) z |= 4'b0100; 
	if(x==?20'b??????1??1??1????0?0) z |= 4'b0010; 
	if(x==?20'b?????????11?1???0??0) z |= 4'b0010; 
	if(x==?20'b?????1???1??1???0??0) z |= 4'b0010; 
	if(x==?20'b?????1????1????1?0?0) z |= 4'b0001; 
	if(x==?20'b?????????11????10??0) z |= 4'b0001; 
	if(x==?20'b??????1???1????10??0) z |= 4'b0001; 
	if(x==?20'b1????1???11????????0) z |= 4'b1000; 
	if(x==?20'b1????11???1????????0) z |= 4'b1000; 
	if(x==?20'b???1??1??11????????0) z |= 4'b0100; 
	if(x==?20'b???1?11??1?????????0) z |= 4'b0100; 
	if(x==?20'b??????1??11?1??????0) z |= 4'b0010; 
	if(x==?20'b?????11??1??1??????0) z |= 4'b0010; 
	if(x==?20'b?????1???11????1???0) z |= 4'b0001; 
	if(x==?20'b?????11???1????1???0) z |= 4'b0001; 
	if(x==?20'b?????11??11?????000?) z |= 4'b1111; 
	if(x==?20'b????????1???????0000) z |= 4'b1000; 
	if(x==?20'b??1?????????????0000) z |= 4'b1000; 
	if(x==?20'b???????????1????0000) z |= 4'b0100; 
	if(x==?20'b?1??????????????0000) z |= 4'b0100; 
	if(x==?20'b??????????????1?0000) z |= 4'b0010; 
	if(x==?20'b????1???????????0000) z |= 4'b0010; 
	if(x==?20'b?????????????1??0000) z |= 4'b0001; 
	if(x==?20'b???????1????????0000) z |= 4'b0001; 
	if(x==?20'b????????1?1??????000) z |= 4'b1000; 
	if(x==?20'b??1???????1??????000) z |= 4'b1000; 
	if(x==?20'b????????11??????0?00) z |= 4'b1000; 
	if(x==?20'b??1???1?????????0?00) z |= 4'b1000; 
	if(x==?20'b?????????1?1?????000) z |= 4'b0100; 
	if(x==?20'b?1???????1???????000) z |= 4'b0100; 
	if(x==?20'b??????????11????0?00) z |= 4'b0100; 
	if(x==?20'b?1???1??????????0?00) z |= 4'b0100; 
	if(x==?20'b??????1???????1??000) z |= 4'b0010; 
	if(x==?20'b????1?1??????????000) z |= 4'b0010; 
	if(x==?20'b??????????1???1?0?00) z |= 4'b0010; 
	if(x==?20'b????11??????????0?00) z |= 4'b0010; 
	if(x==?20'b?????1???????1???000) z |= 4'b0001; 
	if(x==?20'b?????1?1?????????000) z |= 4'b0001; 
	if(x==?20'b?????????1???1??0?00) z |= 4'b0001; 
	if(x==?20'b??????11????????0?00) z |= 4'b0001; 
	if(x==?20'b????????111???????00) z |= 4'b1000; 
	if(x==?20'b??1??????11???????00) z |= 4'b1000; 
	if(x==?20'b??????1?1?1???????00) z |= 4'b1000; 
	if(x==?20'b??1???1???1???????00) z |= 4'b1000; 
	if(x==?20'b?????1??1???????00?0) z |= 4'b1000; 
	if(x==?20'b??1??1??????????00?0) z |= 4'b1000; 
	if(x==?20'b?????????111??????00) z |= 4'b0100; 
	if(x==?20'b?????1???1?1??????00) z |= 4'b0100; 
	if(x==?20'b?1???????11???????00) z |= 4'b0100; 
	if(x==?20'b?1???1???1????????00) z |= 4'b0100; 
	if(x==?20'b??????1????1????00?0) z |= 4'b0100; 
	if(x==?20'b?1????1?????????00?0) z |= 4'b0100; 
	if(x==?20'b??????1???1???1???00) z |= 4'b0010; 
	if(x==?20'b?????11???????1???00) z |= 4'b0010; 
	if(x==?20'b????1?1???1???????00) z |= 4'b0010; 
	if(x==?20'b????111???????????00) z |= 4'b0010; 
	if(x==?20'b?????????1????1?00?0) z |= 4'b0010; 
	if(x==?20'b????1????1??????00?0) z |= 4'b0010; 
	if(x==?20'b?????1???1???1????00) z |= 4'b0001; 
	if(x==?20'b?????11??????1????00) z |= 4'b0001; 
	if(x==?20'b?????1?1?1????????00) z |= 4'b0001; 
	if(x==?20'b?????111??????????00) z |= 4'b0001; 
	if(x==?20'b??????????1??1??00?0) z |= 4'b0001; 
	if(x==?20'b???????1??1?????00?0) z |= 4'b0001; 
	if(x==?20'b????11????1?????0??0) z |= 4'b1000; 
	if(x==?20'b?1???1????1?????0??0) z |= 4'b1000; 
	if(x==?20'b?????1??11??????0??0) z |= 4'b1000; 
	if(x==?20'b??1??1???1??????0??0) z |= 4'b1000; 
	if(x==?20'b?????11?1???????0??0) z |= 4'b1000; 
	if(x==?20'b??1??11?????????0??0) z |= 4'b1000; 
	if(x==?20'b??????1???11????0??0) z |= 4'b0100; 
	if(x==?20'b?????11????1????0??0) z |= 4'b0100; 
	if(x==?20'b?1????1???1?????0??0) z |= 4'b0100; 
	if(x==?20'b??????11?1??????0??0) z |= 4'b0100; 
	if(x==?20'b??1???1??1??????0??0) z |= 4'b0100; 
	if(x==?20'b?1???11?????????0??0) z |= 4'b0100; 
	if(x==?20'b?????????11???1?0??0) z |= 4'b0010; 
	if(x==?20'b?????1???1????1?0??0) z |= 4'b0010; 
	if(x==?20'b??????1??1???1??0??0) z |= 4'b0010; 
	if(x==?20'b????1????11?????0??0) z |= 4'b0010; 
	if(x==?20'b??????1?11??????0??0) z |= 4'b0010; 
	if(x==?20'b????11???1??????0??0) z |= 4'b0010; 
	if(x==?20'b?????1????1???1?0??0) z |= 4'b0001; 
	if(x==?20'b?????????11??1??0??0) z |= 4'b0001; 
	if(x==?20'b??????1???1??1??0??0) z |= 4'b0001; 
	if(x==?20'b?????1????11????0??0) z |= 4'b0001; 
	if(x==?20'b???????1?11?????0??0) z |= 4'b0001; 
	if(x==?20'b??????11??1?????0??0) z |= 4'b0001; 
	if(x==?20'b?????1??111????????0) z |= 4'b1000; 
	if(x==?20'b??1??1???11????????0) z |= 4'b1000; 
	if(x==?20'b?????11?1?1????????0) z |= 4'b1000; 
	if(x==?20'b??1??11???1????????0) z |= 4'b1000; 
	if(x==?20'b??????1??111???????0) z |= 4'b0100; 
	if(x==?20'b?????11??1?1???????0) z |= 4'b0100; 
	if(x==?20'b?1????1??11????????0) z |= 4'b0100; 
	if(x==?20'b?1???11??1?????????0) z |= 4'b0100; 
	if(x==?20'b??????1??11???1????0) z |= 4'b0010; 
	if(x==?20'b?????11??1????1????0) z |= 4'b0010; 
	if(x==?20'b????1?1??11????????0) z |= 4'b0010; 
	if(x==?20'b????111??1?????????0) z |= 4'b0010; 
	if(x==?20'b?????1???11??1?????0) z |= 4'b0001; 
	if(x==?20'b?????11???1??1?????0) z |= 4'b0001; 
	if(x==?20'b?????1?1?11????????0) z |= 4'b0001; 
	if(x==?20'b?????111??1????????0) z |= 4'b0001; 
	if(x==?20'b?11?????????????0?00) z |= 4'b1100; 
	if(x==?20'b????1???1???????0?00) z |= 4'b1010; 
	if(x==?20'b???????1???1????0?00) z |= 4'b0101; 
	if(x==?20'b?????????????11?0?00) z |= 4'b0011; 
	if(x==?20'b??????????1?????0000) z |= 4'b1000; 
	if(x==?20'b?????????1??????0000) z |= 4'b0100; 
	if(x==?20'b??????1?????????0000) z |= 4'b0010; 
	if(x==?20'b?????1??????????0000) z |= 4'b0001; 
	if(x==?20'b?1??1?????????????00) z |= 4'b1000; 
	if(x==?20'b??1????1??????????00) z |= 4'b0100; 
	if(x==?20'b????????1????1????00) z |= 4'b0010; 
	if(x==?20'b???????????1??1???00) z |= 4'b0001; 
	if(x==?20'b?1????????1?????0?00) z |= 4'b1100; 
	if(x==?20'b??1??????1??????0?00) z |= 4'b1100; 
	if(x==?20'b????1?????1?????0?00) z |= 4'b1010; 
	if(x==?20'b??????1?1???????0?00) z |= 4'b1010; 
	if(x==?20'b?????1?????1????0?00) z |= 4'b0101; 
	if(x==?20'b???????1?1??????0?00) z |= 4'b0101; 
	if(x==?20'b?????1????????1?0?00) z |= 4'b0011; 
	if(x==?20'b??????1??????1??0?00) z |= 4'b0011; 
	if(x==?20'b?1??11?????????????0) z |= 4'b1000; 
	if(x==?20'b??1???11???????????0) z |= 4'b0100; 
	if(x==?20'b????????11???1?????0) z |= 4'b0010; 
	if(x==?20'b??????????11??1????0) z |= 4'b0001; 
	if(x==?20'b??1??1????1??????0?0) z |= 4'b1100; 
	if(x==?20'b?1????1??1???????0?0) z |= 4'b1100; 
	if(x==?20'b?????1??1?1??????0?0) z |= 4'b1010; 
	if(x==?20'b????1?1??1???????0?0) z |= 4'b1010; 
	if(x==?20'b??????1??1?1?????0?0) z |= 4'b0101; 
	if(x==?20'b?????1?1??1??????0?0) z |= 4'b0101; 
	if(x==?20'b??????1??1????1??0?0) z |= 4'b0011; 
	if(x==?20'b?????1????1??1???0?0) z |= 4'b0011; 
	if(x==?20'b????1????????????000) z |= 4'b1000; 
	if(x==?20'b?1???????????????000) z |= 4'b1000; 
	if(x==?20'b???????1?????????000) z |= 4'b0100; 
	if(x==?20'b??1??????????????000) z |= 4'b0100; 
	if(x==?20'b?????????????1???000) z |= 4'b0010; 
	if(x==?20'b????????1????????000) z |= 4'b0010; 
	if(x==?20'b??????????????1??000) z |= 4'b0001; 
	if(x==?20'b???????????1?????000) z |= 4'b0001; 
	if(x==?20'b????1????1????????00) z |= 4'b1000; 
	if(x==?20'b?1???????1????????00) z |= 4'b1000; 
	if(x==?20'b????1?1???????????00) z |= 4'b1000; 
	if(x==?20'b?1????1???????????00) z |= 4'b1000; 
	if(x==?20'b???????1??1???????00) z |= 4'b0100; 
	if(x==?20'b??1???????1???????00) z |= 4'b0100; 
	if(x==?20'b?????1?1??????????00) z |= 4'b0100; 
	if(x==?20'b??1??1????????????00) z |= 4'b0100; 
	if(x==?20'b??????????1??1????00) z |= 4'b0010; 
	if(x==?20'b?????1???????1????00) z |= 4'b0010; 
	if(x==?20'b????????1?1???????00) z |= 4'b0010; 
	if(x==?20'b?????1??1?????????00) z |= 4'b0010; 
	if(x==?20'b?????????1????1???00) z |= 4'b0001; 
	if(x==?20'b??????1???????1???00) z |= 4'b0001; 
	if(x==?20'b?????????1?1??????00) z |= 4'b0001; 
	if(x==?20'b??????1????1??????00) z |= 4'b0001; 
	if(x==?20'b?????????11?????0?00) z |= 4'b1100; 
	if(x==?20'b??????1???1?????0?00) z |= 4'b1010; 
	if(x==?20'b?????1???1??????0?00) z |= 4'b0101; 
	if(x==?20'b?????11?????????0?00) z |= 4'b0011; 
	if(x==?20'b????11???????????0?0) z |= 4'b1000; 
	if(x==?20'b?1???1???????????0?0) z |= 4'b1000; 
	if(x==?20'b??????11?????????0?0) z |= 4'b0100; 
	if(x==?20'b??1???1??????????0?0) z |= 4'b0100; 
	if(x==?20'b?????????1???1???0?0) z |= 4'b0010; 
	if(x==?20'b????????11???????0?0) z |= 4'b0010; 
	if(x==?20'b??????????1???1??0?0) z |= 4'b0001; 
	if(x==?20'b??????????11?????0?0) z |= 4'b0001; 
	if(x==?20'b??????1??1??????00?0) z |= 4'b0110; 
	if(x==?20'b?????1????1?????00?0) z |= 4'b1001; 
	if(x==?20'b????11???1?????????0) z |= 4'b1000; 
	if(x==?20'b?1???1???1?????????0) z |= 4'b1000; 
	if(x==?20'b????111????????????0) z |= 4'b1000; 
	if(x==?20'b?1???11????????????0) z |= 4'b1000; 
	if(x==?20'b??????11??1????????0) z |= 4'b0100; 
	if(x==?20'b??1???1???1????????0) z |= 4'b0100; 
	if(x==?20'b?????111???????????0) z |= 4'b0100; 
	if(x==?20'b??1??11????????????0) z |= 4'b0100; 
	if(x==?20'b?????????11??1?????0) z |= 4'b0010; 
	if(x==?20'b?????1???1???1?????0) z |= 4'b0010; 
	if(x==?20'b????????111????????0) z |= 4'b0010; 
	if(x==?20'b?????1??11?????????0) z |= 4'b0010; 
	if(x==?20'b?????????11???1????0) z |= 4'b0001; 
	if(x==?20'b??????1???1???1????0) z |= 4'b0001; 
	if(x==?20'b?????????111???????0) z |= 4'b0001; 
	if(x==?20'b??????1???11???????0) z |= 4'b0001; 
	if(x==?20'b??????1??11?????0??0) z |= 4'b0110; 
	if(x==?20'b?????11??1??????0??0) z |= 4'b0110; 
	if(x==?20'b?????1???11?????0??0) z |= 4'b1001; 
	if(x==?20'b?????11???1?????0??0) z |= 4'b1001; 
	if(x==?20'b?????11??1?????????0) z |= 4'b1000; 
	if(x==?20'b?????11???1????????0) z |= 4'b0100; 
	if(x==?20'b?????1???11????????0) z |= 4'b0010; 
	if(x==?20'b??????1??11????????0) z |= 4'b0001; 
	if(x==?20'b??????????1??????000) z |= 4'b0110; 
	if(x==?20'b?????1???????????000) z |= 4'b0110; 
	if(x==?20'b?????????1???????000) z |= 4'b1001; 
	if(x==?20'b??????1??????????000) z |= 4'b1001; 
	if(x==?20'b?????1????1???????00) z |= 4'b0110; 
	if(x==?20'b??????1??1????????00) z |= 4'b1001; 
	if(x==?20'b?????11??????????0?0) z |= 4'b1100; 
	if(x==?20'b?????1???1???????0?0) z |= 4'b1010; 
	if(x==?20'b??????1???1??????0?0) z |= 4'b0101; 
	if(x==?20'b?????????11??????0?0) z |= 4'b0011; 
	if(x==?20'b?????1????????????00) z |= 4'b1000; 
	if(x==?20'b??????1???????????00) z |= 4'b0100; 
	if(x==?20'b?????????1????????00) z |= 4'b0010; 
	if(x==?20'b??????????1???????00) z |= 4'b0001; 
end 
endmodule