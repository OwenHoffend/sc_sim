module gb4_opt_pairs(
    input [19:0] x,
    output logic [3:0] z
);
always_comb begin 
	 z = 4'b0000;
	if(x==?20'b1???1?00100??1110011) z |= 4'b1000; 
	if(x==?20'b???100?1?001111?0011) z |= 4'b0100; 
	if(x==?20'b?111110?110?011?1?00) z |= 4'b0100; 
	if(x==?20'b111??011?011?1101?00) z |= 4'b1000; 
	if(x==?20'b??1?00?1111?111?0010) z |= 4'b0100; 
	if(x==?20'b?1??1?00?111?1110010) z |= 4'b1000; 
	if(x==?20'b?111110?110?110?1?00) z |= 4'b0100; 
	if(x==?20'b111??011?011?0111?00) z |= 4'b1000; 
	if(x==?20'b??1?1?00100??1110011) z |= 4'b1000; 
	if(x==?20'b?1??00?1?001111?0011) z |= 4'b0100; 
	if(x==?20'b?????0111110?1101000) z |= 4'b1000; 
	if(x==?20'b????110?0111011?1000) z |= 4'b0100; 
	if(x==?20'b????110?0111110?1000) z |= 4'b0100; 
	if(x==?20'b?????0111110?0111000) z |= 4'b1000; 
	if(x==?20'b?1?1001?111?111?0?10) z |= 4'b0100; 
	if(x==?20'b1?1??100?111?1110?10) z |= 4'b1000; 
	if(x==?20'b????00?1000?111?0011) z |= 4'b0100; 
	if(x==?20'b????1?00?000?1110011) z |= 4'b1000; 
	if(x==?20'b???1?0?1000?111?0011) z |= 4'b0100; 
	if(x==?20'b1???1?0??000?1110011) z |= 4'b1000; 
	if(x==?20'b?1?110??100?001?1100) z |= 4'b0100; 
	if(x==?20'b1?1???01?001?1001100) z |= 4'b1000; 
	if(x==?20'b?????0?10001111?0011) z |= 4'b0100; 
	if(x==?20'b????1?0?1000?1110011) z |= 4'b1000; 
	if(x==?20'b???10???0001111?0011) z |= 4'b0100; 
	if(x==?20'b1??????01000?1110011) z |= 4'b1000; 
	if(x==?20'b?1?110??100?100?1100) z |= 4'b0100; 
	if(x==?20'b1?1???01?001?0011100) z |= 4'b1000; 
	if(x==?20'b????0??10001111?0011) z |= 4'b0100; 
	if(x==?20'b????1??01000?1110011) z |= 4'b1000; 
	if(x==?20'b?1???0?1000?111?0011) z |= 4'b0100; 
	if(x==?20'b??1?1?0??000?1110011) z |= 4'b1000; 
	if(x==?20'b???1???10001111?0011) z |= 4'b0100; 
	if(x==?20'b1???1???1000?1110011) z |= 4'b1000; 
	if(x==?20'b?1?1001?110111??1?10) z |= 4'b0100; 
	if(x==?20'b?11100??110?011?101?) z |= 4'b0100; 
	if(x==?20'b111???00?011?110101?) z |= 4'b1000; 
	if(x==?20'b?11100??011?011?101?) z |= 4'b0100; 
	if(x==?20'b111???00?110?110101?) z |= 4'b1000; 
	if(x==?20'b????010?011101??0100) z |= 4'b0100; 
	if(x==?20'b?????0101110??100100) z |= 4'b1000; 
	if(x==?20'b?1??0???0001111?0011) z |= 4'b0100; 
	if(x==?20'b??1????01000?1110011) z |= 4'b1000; 
	if(x==?20'b?11100??110?110?101?) z |= 4'b0100; 
	if(x==?20'b111???00?011?011101?) z |= 4'b1000; 
	if(x==?20'b1?1??1001011?11?1?10) z |= 4'b1000; 
	if(x==?20'b?11100??011?110?101?) z |= 4'b0100; 
	if(x==?20'b?1?1001?11?1011?1?10) z |= 4'b0100; 
	if(x==?20'b?????01?1110?1010100) z |= 4'b1000; 
	if(x==?20'b???100?1111?00??0001) z |= 4'b0100; 
	if(x==?20'b1???1000?011??111?10) z |= 4'b1000; 
	if(x==?20'b???1001??001111?0?11) z |= 4'b0100; 
	if(x==?20'b?????10?0111101?0100) z |= 4'b0100; 
	if(x==?20'b1???1?00?111??000001) z |= 4'b1000; 
	if(x==?20'b111???00?110?011101?) z |= 4'b1000; 
	if(x==?20'b1????100100??1110?11) z |= 4'b1000; 
	if(x==?20'b111???001110?11?101?) z |= 4'b1000; 
	if(x==?20'b?11100??0111?11?101?) z |= 4'b0100; 
	if(x==?20'b111???0?1110?110101?) z |= 4'b1000; 
	if(x==?20'b?1?????10001111?0011) z |= 4'b0100; 
	if(x==?20'b?111?0??0111011?101?) z |= 4'b0100; 
	if(x==?20'b??1?1???1000?1110011) z |= 4'b1000; 
	if(x==?20'b??????101101?1010100) z |= 4'b1000; 
	if(x==?20'b????01??1011101?0100) z |= 4'b0100; 
	if(x==?20'b???10001110??11?1?10) z |= 4'b0100; 
	if(x==?20'b?????0001110?110101?) z |= 4'b1000; 
	if(x==?20'b1?1??1001?11?0111?10) z |= 4'b1000; 
	if(x==?20'b????000?0111011?101?) z |= 4'b0100; 
	if(x==?20'b????010?0111?10?0100) z |= 4'b0100; 
	if(x==?20'b?????0101110?01?0100) z |= 4'b1000; 
	if(x==?20'b?11??001?001??011100) z |= 4'b1100; 
	if(x==?20'b?111?0??0111110?101?) z |= 4'b0100; 
	if(x==?20'b?????10?0111010?0100) z |= 4'b0100; 
	if(x==?20'b1???1000??11?1101?10) z |= 4'b1000; 
	if(x==?20'b?????01?1110?0100100) z |= 4'b1000; 
	if(x==?20'b????100?011101??1100) z |= 4'b0100; 
	if(x==?20'b111???0?1110?011101?) z |= 4'b1000; 
	if(x==?20'b?????0011110??101100) z |= 4'b1000; 
	if(x==?20'b????00?1111?000?0001) z |= 4'b0100; 
	if(x==?20'b????1?00?111?0000001) z |= 4'b1000; 
	if(x==?20'b111????01110?110101?) z |= 4'b1000; 
	if(x==?20'b?????001110??0101100) z |= 4'b1000; 
	if(x==?20'b?1110???0111011?101?) z |= 4'b0100; 
	if(x==?20'b????100??011010?1100) z |= 4'b0100; 
	if(x==?20'b??1?001?111?111?0?10) z |= 4'b0100; 
	if(x==?20'b????000?0111110?101?) z |= 4'b0100; 
	if(x==?20'b???1000111??110?1?10) z |= 4'b0100; 
	if(x==?20'b?????0001110?011101?) z |= 4'b1000; 
	if(x==?20'b???100?1111??00?0001) z |= 4'b0100; 
	if(x==?20'b????01??1011010?0100) z |= 4'b0100; 
	if(x==?20'b??1?0001110?11??1?10) z |= 4'b0100; 
	if(x==?20'b?1??0001110?11??1?10) z |= 4'b0100; 
	if(x==?20'b??????101101?0100100) z |= 4'b1000; 
	if(x==?20'b?1???100?111?1110?10) z |= 4'b1000; 
	if(x==?20'b1???1?00?111?00?0001) z |= 4'b1000; 
	if(x==?20'b?11?100?100??01?1100) z |= 4'b1100; 
	if(x==?20'b???1?0?1111?000?0001) z |= 4'b0100; 
	if(x==?20'b????100?01111?0?1100) z |= 4'b0100; 
	if(x==?20'b1???1?0??111?0000001) z |= 4'b1000; 
	if(x==?20'b?????0011110?0?11100) z |= 4'b1000; 
	if(x==?20'b?1??00?1111?00??0001) z |= 4'b0100; 
	if(x==?20'b?1??1000?011??111?10) z |= 4'b1000; 
	if(x==?20'b?1??001??001111?0?11) z |= 4'b0100; 
	if(x==?20'b??1?1?00?111??000001) z |= 4'b1000; 
	if(x==?20'b?1110???0111110?101?) z |= 4'b0100; 
	if(x==?20'b??1??100100??1110?11) z |= 4'b1000; 
	if(x==?20'b111????01110?011101?) z |= 4'b1000; 
	if(x==?20'b??1101??010?101??100) z |= 4'b0100; 
	if(x==?20'b11????10?010?101?100) z |= 4'b1000; 
	if(x==?20'b1?1?1??0100??1110?11) z |= 4'b1000; 
	if(x==?20'b1?????001110?110101?) z |= 4'b1000; 
	if(x==?20'b?1?10??1?001111?0?11) z |= 4'b0100; 
	if(x==?20'b?1?1?01??001111?0?11) z |= 4'b0100; 
	if(x==?20'b1?1??10?100??1110?11) z |= 4'b1000; 
	if(x==?20'b?1?1001?0??1111?0?11) z |= 4'b0100; 
	if(x==?20'b1?1??1001??0?1110?11) z |= 4'b1000; 
	if(x==?20'b?11??001?001?10011?0) z |= 4'b1100; 
	if(x==?20'b??1100??010?101?011?) z |= 4'b0100; 
	if(x==?20'b??1?1000?011?11?1?10) z |= 4'b1000; 
	if(x==?20'b???10??1111?000?0001) z |= 4'b0100; 
	if(x==?20'b11????00?010?101011?) z |= 4'b1000; 
	if(x==?20'b1???1??0?111?0000001) z |= 4'b1000; 
	if(x==?20'b??1?000111??011?1?10) z |= 4'b0100; 
	if(x==?20'b?1??000111??011?1?10) z |= 4'b0100; 
	if(x==?20'b?111010??10?01???100) z |= 4'b0100; 
	if(x==?20'b?1??1000??11?1101?10) z |= 4'b1000; 
	if(x==?20'b1?????001110?011101?) z |= 4'b1000; 
	if(x==?20'b111??010?01???10?100) z |= 4'b1000; 
	if(x==?20'b??1?10??100?001?1100) z |= 4'b0100; 
	if(x==?20'b?1????01?001?1001100) z |= 4'b1000; 
	if(x==?20'b??1101??010?010??100) z |= 4'b0100; 
	if(x==?20'b?1110??11101011?1?1?) z |= 4'b0100; 
	if(x==?20'b111?1??01011?1101?1?) z |= 4'b1000; 
	if(x==?20'b11????10?010?010?100) z |= 4'b1000; 
	if(x==?20'b?1??00?1111??00?0001) z |= 4'b0100; 
	if(x==?20'b??1?1?00?111?00?0001) z |= 4'b1000; 
	if(x==?20'b??1110??10??010?1100) z |= 4'b0100; 
	if(x==?20'b??1100??010?010?011?) z |= 4'b0100; 
	if(x==?20'b?1???0?1111?000?0001) z |= 4'b0100; 
	if(x==?20'b?111?10??10?101??100) z |= 4'b0100; 
	if(x==?20'b??1?1?0??111?0000001) z |= 4'b1000; 
	if(x==?20'b??1?10??100?100?1100) z |= 4'b0100; 
	if(x==?20'b111??01??01??101?100) z |= 4'b1000; 
	if(x==?20'b??1?1000??11?0111?10) z |= 4'b1000; 
	if(x==?20'b11????01??01?0101100) z |= 4'b1000; 
	if(x==?20'b11????00?010?010011?) z |= 4'b1000; 
	if(x==?20'b?1110??11101110?1?1?) z |= 4'b0100; 
	if(x==?20'b??1100??101?101?011?) z |= 4'b0100; 
	if(x==?20'b?1????01?001?0011100) z |= 4'b1000; 
	if(x==?20'b11????00?101?101011?) z |= 4'b1000; 
	if(x==?20'b??11?011111?111???10) z |= 4'b0100; 
	if(x==?20'b?11?01??010?101??100) z |= 4'b0100; 
	if(x==?20'b111?1??01011?0111?1?) z |= 4'b1000; 
	if(x==?20'b???10??100??111?0011) z |= 4'b0100; 
	if(x==?20'b?11???10?010?101?100) z |= 4'b1000; 
	if(x==?20'b??11111?0?01111???01) z |= 4'b0100; 
	if(x==?20'b??1???001110?110101?) z |= 4'b1000; 
	if(x==?20'b1???1??0??00?1110011) z |= 4'b1000; 
	if(x==?20'b11??110??111?111??10) z |= 4'b1000; 
	if(x==?20'b11???11110?0?111??01) z |= 4'b1000; 
	if(x==?20'b?11100??010?01??011?) z |= 4'b0100; 
	if(x==?20'b111???00?010??10011?) z |= 4'b1000; 
	if(x==?20'b?111010??10??10??100) z |= 4'b0100; 
	if(x==?20'b?11?00??010?101?011?) z |= 4'b0100; 
	if(x==?20'b?1??0??1111?000?0001) z |= 4'b0100; 
	if(x==?20'b111??010?01??01??100) z |= 4'b1000; 
	if(x==?20'b?11???00?010?101011?) z |= 4'b1000; 
	if(x==?20'b??1?1??0?111?0000001) z |= 4'b1000; 
	if(x==?20'b?111?10??10?010??100) z |= 4'b0100; 
	if(x==?20'b111??01??01??010?100) z |= 4'b1000; 
	if(x==?20'b?1?1001?111?0?0?0?01) z |= 4'b0100; 
	if(x==?20'b??1100??101?010?011?) z |= 4'b0100; 
	if(x==?20'b1?1??100?111?0?00?01) z |= 4'b1000; 
	if(x==?20'b??1???001110?011101?) z |= 4'b1000; 
	if(x==?20'b11????00?101?010011?) z |= 4'b1000; 
	if(x==?20'b11????0?1101?101011?) z |= 4'b1000; 
	if(x==?20'b?11?01??010?010??100) z |= 4'b0100; 
	if(x==?20'b?111?0??010?101?011?) z |= 4'b0100; 
	if(x==?20'b??11?0??1011101?011?) z |= 4'b0100; 
	if(x==?20'b?11100???10?101?011?) z |= 4'b0100; 
	if(x==?20'b111???0??010?101011?) z |= 4'b1000; 
	if(x==?20'b?11100??01??101?011?) z |= 4'b0100; 
	if(x==?20'b?11???10?010?010?100) z |= 4'b1000; 
	if(x==?20'b111???00?01??101011?) z |= 4'b1000; 
	if(x==?20'b111???00??10?101011?) z |= 4'b1000; 
	if(x==?20'b????1101?010?1?1010?) z |= 4'b1000; 
	if(x==?20'b?11?10??10??010?1100) z |= 4'b0100; 
	if(x==?20'b?11100??101?01??011?) z |= 4'b0100; 
	if(x==?20'b?11?00??010?010?011?) z |= 4'b0100; 
	if(x==?20'b?11100??01?101??011?) z |= 4'b0100; 
	if(x==?20'b111???00?101??10011?) z |= 4'b1000; 
	if(x==?20'b111???001?10??10011?) z |= 4'b1000; 
	if(x==?20'b?11???01??01?0101100) z |= 4'b1000; 
	if(x==?20'b?11???00?010?010011?) z |= 4'b1000; 
	if(x==?20'b?11?00??101?101?011?) z |= 4'b0100; 
	if(x==?20'b?11???00?101?101011?) z |= 4'b1000; 
	if(x==?20'b?1?111?1?00111??1?01) z |= 4'b0100; 
	if(x==?20'b??1?001?1101?11?1?10) z |= 4'b0100; 
	if(x==?20'b?11100??010??10?011?) z |= 4'b0100; 
	if(x==?20'b?1???1001011?11?1?10) z |= 4'b1000; 
	if(x==?20'b?11??011111?111???10) z |= 4'b0100; 
	if(x==?20'b1?1?1?11100???111?01) z |= 4'b1000; 
	if(x==?20'b?1??0??100??111?0011) z |= 4'b0100; 
	if(x==?20'b?11?111?0?01111???01) z |= 4'b0100; 
	if(x==?20'b?111?0??010?010?011?) z |= 4'b0100; 
	if(x==?20'b??11?0??1011010?011?) z |= 4'b0100; 
	if(x==?20'b??1?1??0??00?1110011) z |= 4'b1000; 
	if(x==?20'b111???00?010?01?011?) z |= 4'b1000; 
	if(x==?20'b?11?110??111?111??10) z |= 4'b1000; 
	if(x==?20'b11????0?1101?010011?) z |= 4'b1000; 
	if(x==?20'b?11??11110?0?111??01) z |= 4'b1000; 
	if(x==?20'b?????01?0001111?0?11) z |= 4'b0100; 
	if(x==?20'b?11100???10?010?011?) z |= 4'b0100; 
	if(x==?20'b?11100??01??010?011?) z |= 4'b0100; 
	if(x==?20'b?????10?1000?1110?11) z |= 4'b1000; 
	if(x==?20'b111???0??010?010011?) z |= 4'b1000; 
	if(x==?20'b111???00?01??010011?) z |= 4'b1000; 
	if(x==?20'b?111?0??101?101?011?) z |= 4'b0100; 
	if(x==?20'b111???0??101?101011?) z |= 4'b1000; 
	if(x==?20'b111???00??10?010011?) z |= 4'b1000; 
	if(x==?20'b111???0?1?10?101011?) z |= 4'b1000; 
	if(x==?20'b?111?0??01?1101?011?) z |= 4'b0100; 
	if(x==?20'b?111?0??101101??011?) z |= 4'b0100; 
	if(x==?20'b1?1?1?11100??11?1?01) z |= 4'b1000; 
	if(x==?20'b??1?001?11?1110?1?10) z |= 4'b0100; 
	if(x==?20'b111???0?1101??10011?) z |= 4'b1000; 
	if(x==?20'b?11?00??101?010?011?) z |= 4'b0100; 
	if(x==?20'b?1?111?1?001?11?1?01) z |= 4'b0100; 
	if(x==?20'b?11???00?101?010011?) z |= 4'b1000; 
	if(x==?20'b?11???0?1101?101011?) z |= 4'b1000; 
	if(x==?20'b?11??0??1011101?011?) z |= 4'b0100; 
	if(x==?20'b?????001110???011100) z |= 4'b1000; 
	if(x==?20'b?1???1001?11?0111?10) z |= 4'b1000; 
	if(x==?20'b?????00111?0??011100) z |= 4'b1000; 
	if(x==?20'b???10001?1??101??110) z |= 4'b0100; 
	if(x==?20'b1???1000??1??101?110) z |= 4'b1000; 
	if(x==?20'b?11100??101??10?011?) z |= 4'b0100; 
	if(x==?20'b?11100??01?1?10?011?) z |= 4'b0100; 
	if(x==?20'b111???00?101?01?011?) z |= 4'b1000; 
	if(x==?20'b111???001?10?01?011?) z |= 4'b1000; 
	if(x==?20'b??1?0???0001111?0?11) z |= 4'b0100; 
	if(x==?20'b?111?0??101?010?011?) z |= 4'b0100; 
	if(x==?20'b?111?0??01?1010?011?) z |= 4'b0100; 
	if(x==?20'b?1?????01000?1110?11) z |= 4'b1000; 
	if(x==?20'b111???0??101?010011?) z |= 4'b1000; 
	if(x==?20'b111???0?1?10?010011?) z |= 4'b1000; 
	if(x==?20'b???10??11101000?1?01) z |= 4'b0100; 
	if(x==?20'b1???1??01011?0001?01) z |= 4'b1000; 
	if(x==?20'b?111?0?1110?011?1?1?) z |= 4'b0100; 
	if(x==?20'b?11111??011?011?1?0?) z |= 4'b0100; 
	if(x==?20'b????10??001?001?1100) z |= 4'b0100; 
	if(x==?20'b111???11?110?1101?0?) z |= 4'b1000; 
	if(x==?20'b??????01?100?1001100) z |= 4'b1001; 
	if(x==?20'b1?1?1??01110?1101?1?) z |= 4'b1000; 
	if(x==?20'b111?1?0??011?1101?1?) z |= 4'b1000; 
	if(x==?20'b?1?10??10111011?1?1?) z |= 4'b0100; 
	if(x==?20'b????100?0?11?01?1100) z |= 4'b0100; 
	if(x==?20'b?11??0??1011010?011?) z |= 4'b0100; 
	if(x==?20'b????100??011?01?1100) z |= 4'b0100; 
	if(x==?20'b?11???0?1101?010011?) z |= 4'b1000; 
	if(x==?20'b111???111110??111?0?) z |= 4'b1000; 
	if(x==?20'b?1?1001??0??111?0?11) z |= 4'b0100; 
	if(x==?20'b???10001?1??010??110) z |= 4'b0100; 
	if(x==?20'b?1?10??1110100??1?01) z |= 4'b0100; 
	if(x==?20'b1?1??100??0??1110?11) z |= 4'b1000; 
	if(x==?20'b1?1?1??01011??001?01) z |= 4'b1000; 
	if(x==?20'b1???1000??1??010?110) z |= 4'b1000; 
	if(x==?20'b?11111?111010?0?1?1?) z |= 4'b0100; 
	if(x==?20'b?111?0?1011?011?1?1?) z |= 4'b0100; 
	if(x==?20'b111?1?0??110?1101?1?) z |= 4'b1000; 
	if(x==?20'b111?1?111011?0?01?1?) z |= 4'b1000; 
	if(x==?20'b?111?0??1011?10?011?) z |= 4'b0100; 
	if(x==?20'b111???0?1101?01?011?) z |= 4'b1000; 
	if(x==?20'b?111?0?1110?110?1?1?) z |= 4'b0100; 
	if(x==?20'b?1??1??0100??1110?11) z |= 4'b1000; 
	if(x==?20'b1???1?00?000??111?11) z |= 4'b1000; 
	if(x==?20'b??1?0??1?001111?0?11) z |= 4'b0100; 
	if(x==?20'b?11111??011?110?1?0?) z |= 4'b0100; 
	if(x==?20'b??????01?100?0011100) z |= 4'b1000; 
	if(x==?20'b?1?10??10111110?1?1?) z |= 4'b0100; 
	if(x==?20'b????10??001?100?1100) z |= 4'b0110; 
	if(x==?20'b??1??01??001111?0?11) z |= 4'b0100; 
	if(x==?20'b?1???10?100??1110?11) z |= 4'b1000; 
	if(x==?20'b111???11?110?0111?0?) z |= 4'b1000; 
	if(x==?20'b1?1?1??01110?0111?1?) z |= 4'b1000; 
	if(x==?20'b111?1?0??011?0111?1?) z |= 4'b1000; 
	if(x==?20'b??1?001?0??1111?0?11) z |= 4'b0100; 
	if(x==?20'b?1???1001??0?1110?11) z |= 4'b1000; 
	if(x==?20'b??????001101?101011?) z |= 4'b1000; 
	if(x==?20'b?11111??0111?11?1?0?) z |= 4'b0100; 
	if(x==?20'b?111?0?1011?110?1?1?) z |= 4'b0100; 
	if(x==?20'b????00?1000?011?1?11) z |= 4'b0100; 
	if(x==?20'b????00??1011101?011?) z |= 4'b0100; 
	if(x==?20'b????1?00?000?1101?11) z |= 4'b1000; 
	if(x==?20'b????1110?011??11100?) z |= 4'b1000; 
	if(x==?20'b??????01110??1001100) z |= 4'b1000; 
	if(x==?20'b??????0111?0?1001100) z |= 4'b1000; 
	if(x==?20'b?1??0001?1??101??110) z |= 4'b0100; 
	if(x==?20'b??1?1000??1??101?110) z |= 4'b1000; 
	if(x==?20'b111?1?0??110?0111?1?) z |= 4'b1000; 
	if(x==?20'b????10??0?11001?1100) z |= 4'b0100; 
	if(x==?20'b????10???011001?1100) z |= 4'b0100; 
	if(x==?20'b???1001?111?00??0?01) z |= 4'b0100; 
	if(x==?20'b111?1?0?1110?11?1?1?) z |= 4'b1000; 
	if(x==?20'b???100?1000??11?1?11) z |= 4'b0100; 
	if(x==?20'b?1110??1011?011?1?1?) z |= 4'b0100; 
	if(x==?20'b111?1??0?110?1101?1?) z |= 4'b1000; 
	if(x==?20'b??????001110?101011?) z |= 4'b1000; 
	if(x==?20'b1????100?111??000?01) z |= 4'b1000; 
	if(x==?20'b?111?0?10111?11?1?1?) z |= 4'b0100; 
	if(x==?20'b????00??0111101?011?) z |= 4'b0100; 
	if(x==?20'b?1?10?1?11010?0?1?01) z |= 4'b0100; 
	if(x==?20'b???1?0?1000?011?1?11) z |= 4'b0100; 
	if(x==?20'b1???1?0??000?1101?11) z |= 4'b1000; 
	if(x==?20'b1?1??1?01011?0?01?01) z |= 4'b1000; 
	if(x==?20'b?1??0??11101000?1?01) z |= 4'b0100; 
	if(x==?20'b??1?1??01011?0001?01) z |= 4'b1000; 
	if(x==?20'b11????01??01??011100) z |= 4'b1000; 
	if(x==?20'b????00?1000?110?1?11) z |= 4'b0100; 
	if(x==?20'b????0111110??11?100?) z |= 4'b0100; 
	if(x==?20'b?????1011110?10101??) z |= 4'b1000; 
	if(x==?20'b????101?0111101?01??) z |= 4'b0100; 
	if(x==?20'b????1?00?000?0111?11) z |= 4'b1000; 
	if(x==?20'b??????01110??0011100) z |= 4'b1000; 
	if(x==?20'b?????111110?011?100?) z |= 4'b0100; 
	if(x==?20'b????10??0?11100?1100) z |= 4'b0100; 
	if(x==?20'b????10???011100?1100) z |= 4'b0100; 
	if(x==?20'b?1?10??11101?00?1?01) z |= 4'b0100; 
	if(x==?20'b??????0111?0?0011100) z |= 4'b1000; 
	if(x==?20'b1?1?1??01011?00?1?01) z |= 4'b1000; 
	if(x==?20'b?1110??1011?110?1?1?) z |= 4'b0100; 
	if(x==?20'b????111??011?110100?) z |= 4'b1000; 
	if(x==?20'b????00??1011010?011?) z |= 4'b0100; 
	if(x==?20'b??????001101?010011?) z |= 4'b1000; 
	if(x==?20'b?1?1???11101000?1?01) z |= 4'b0100; 
	if(x==?20'b1?1?1???1011?0001?01) z |= 4'b1000; 
	if(x==?20'b???1?0?1000?110?1?11) z |= 4'b0100; 
	if(x==?20'b?1??0001?1??010??110) z |= 4'b0100; 
	if(x==?20'b111?1??0?110?0111?1?) z |= 4'b1000; 
	if(x==?20'b??1?1000??1??010?110) z |= 4'b1000; 
	if(x==?20'b111?1??01110?11?1?1?) z |= 4'b1000; 
	if(x==?20'b111?1?111??0?1101??1) z |= 4'b1000; 
	if(x==?20'b1???1?0??000?0111?11) z |= 4'b1000; 
	if(x==?20'b?1110??10111?11?1?1?) z |= 4'b0100; 
	if(x==?20'b?11111?10??1011?1??1) z |= 4'b0100; 
	if(x==?20'b????00??0111010?011?) z |= 4'b0100; 
	if(x==?20'b??1110??10???01?1100) z |= 4'b0100; 
	if(x==?20'b??????001110?010011?) z |= 4'b1000; 
	if(x==?20'b???100?1110?00??1?01) z |= 4'b0100; 
	if(x==?20'b111?1???1110?1101?1?) z |= 4'b1000; 
	if(x==?20'b?????111110?110?100?) z |= 4'b0100; 
	if(x==?20'b?111???10111011?1?1?) z |= 4'b0100; 
	if(x==?20'b????001?111?000?0?01) z |= 4'b0100; 
	if(x==?20'b1???1?00?011??001?01) z |= 4'b1000; 
	if(x==?20'b?????100?111?0000?01) z |= 4'b1000; 
	if(x==?20'b?111?1??010?01???100) z |= 4'b0100; 
	if(x==?20'b?11101??01??01???100) z |= 4'b0100; 
	if(x==?20'b1???1?001?0??1101?11) z |= 4'b1000; 
	if(x==?20'b????111??011?011100?) z |= 4'b1000; 
	if(x==?20'b111???1??010??10?100) z |= 4'b1000; 
	if(x==?20'b???1001?111??00?0?01) z |= 4'b0100; 
	if(x==?20'b???100?1?0?1011?1?11) z |= 4'b0100; 
	if(x==?20'b111???10??10??10?100) z |= 4'b1000; 
	if(x==?20'b1????100?111?00?0?01) z |= 4'b1000; 
	if(x==?20'b??1100??1011?1??011?) z |= 4'b0100; 
	if(x==?20'b?11111?10??1110?1??1) z |= 4'b0100; 
	if(x==?20'b???1?01?111?000?0?01) z |= 4'b0100; 
	if(x==?20'b11????001101??1?011?) z |= 4'b1000; 
	if(x==?20'b?1?1111??0?1111???01) z |= 4'b0100; 
	if(x==?20'b1?1??1111?0??111??01) z |= 4'b1000; 
	if(x==?20'b111?1?111??0?0111??1) z |= 4'b1000; 
	if(x==?20'b1????10??111?0000?01) z |= 4'b1000; 
	if(x==?20'b?????1101110?11010??) z |= 4'b1000; 
	if(x==?20'b?111???10111110?1?1?) z |= 4'b0100; 
	if(x==?20'b????011?0111011?10??) z |= 4'b0100; 
	if(x==?20'b?1??001?111?00??0?01) z |= 4'b0100; 
	if(x==?20'b??1?001?111?0?0?0?01) z |= 4'b0100; 
	if(x==?20'b?111??1?1101011?1?1?) z |= 4'b0100; 
	if(x==?20'b?1??00?1000??11?1?11) z |= 4'b0100; 
	if(x==?20'b??1?1?00?000?11?1?11) z |= 4'b1000; 
	if(x==?20'b111?1???1110?0111?1?) z |= 4'b1000; 
	if(x==?20'b?1???100?111?0?00?01) z |= 4'b1000; 
	if(x==?20'b??1??100?111??000?01) z |= 4'b1000; 
	if(x==?20'b111??1??1011?1101?1?) z |= 4'b1000; 
	if(x==?20'b??????001101?00001?1) z |= 4'b1000; 
	if(x==?20'b1???1?0?1110?1101?1?) z |= 4'b1000; 
	if(x==?20'b?1???0?1000?011?1?11) z |= 4'b0100; 
	if(x==?20'b??1?1?0??000?1101?11) z |= 4'b1000; 
	if(x==?20'b11????10?101?101?10?) z |= 4'b1000; 
	if(x==?20'b????00??1011000?01?1) z |= 4'b0100; 
	if(x==?20'b??1101??101?101??10?) z |= 4'b0100; 
	if(x==?20'b???1?0?10111011?1?1?) z |= 4'b0100; 
	if(x==?20'b?1?10??1111?00??0?01) z |= 4'b0100; 
	if(x==?20'b???100?1?0?1110?1?11) z |= 4'b0100; 
	if(x==?20'b?1?1001?111??0??0?01) z |= 4'b0100; 
	if(x==?20'b?111?1??01??101??100) z |= 4'b0100; 
	if(x==?20'b1?1?1??0?111??000?01) z |= 4'b1000; 
	if(x==?20'b?1?111?111?100??1?10) z |= 4'b0100; 
	if(x==?20'b111???1???10?101?100) z |= 4'b1000; 
	if(x==?20'b1???1?001?0??0111?11) z |= 4'b1000; 
	if(x==?20'b1?1?1?111?11??001?10) z |= 4'b1000; 
	if(x==?20'b1?1??100?111??0?0?01) z |= 4'b1000; 
	if(x==?20'b?1?1?01?111?00??0?01) z |= 4'b0100; 
	if(x==?20'b??????001110?00010?1) z |= 4'b1000; 
	if(x==?20'b????00?1110?000?1?01) z |= 4'b0100; 
	if(x==?20'b????00??0111000?10?1) z |= 4'b0100; 
	if(x==?20'b1?1??10??111??000?01) z |= 4'b1000; 
	if(x==?20'b????011?0111110?10??) z |= 4'b0100; 
	if(x==?20'b????1?00?011?0001?01) z |= 4'b1000; 
	if(x==?20'b?111??1?1101110?1?1?) z |= 4'b0100; 
	if(x==?20'b????001?00??111?0?11) z |= 4'b0100; 
	if(x==?20'b?????1101110?01110??) z |= 4'b1000; 
	if(x==?20'b?????100??00?1110?11) z |= 4'b1000; 
	if(x==?20'b?1???0?1000?110?1?11) z |= 4'b0100; 
	if(x==?20'b???100?1110??00?1?01) z |= 4'b0100; 
	if(x==?20'b???1?0?10111110?1?1?) z |= 4'b0100; 
	if(x==?20'b111??1??1011?0111?1?) z |= 4'b1000; 
	if(x==?20'b1???1?00?011?00?1?01) z |= 4'b1000; 
	if(x==?20'b?1111???10??0?1?1100) z |= 4'b0100; 
	if(x==?20'b??1?11?1?00111??1?01) z |= 4'b0100; 
	if(x==?20'b1???1?0?1110?0111?1?) z |= 4'b1000; 
	if(x==?20'b????1110111??11010??) z |= 4'b1000; 
	if(x==?20'b???1?0?1110?000?1?01) z |= 4'b0100; 
	if(x==?20'b?111?1??010??10??100) z |= 4'b0100; 
	if(x==?20'b??1?1?0??000?0111?11) z |= 4'b1000; 
	if(x==?20'b111????1??01??101100) z |= 4'b1000; 
	if(x==?20'b?1??1?11100???111?01) z |= 4'b1000; 
	if(x==?20'b????0111?111011?10??) z |= 4'b0100; 
	if(x==?20'b1???1?0??011?0001?01) z |= 4'b1000; 
	if(x==?20'b??1?00?1110?00??1?01) z |= 4'b0100; 
	if(x==?20'b?1??00?1110?00??1?01) z |= 4'b0100; 
	if(x==?20'b111???1??010?01??100) z |= 4'b1000; 
	if(x==?20'b1???1?00??11?0001?01) z |= 4'b1000; 
	if(x==?20'b??1101??101?010??10?) z |= 4'b0100; 
	if(x==?20'b???1?01?00??111?0?11) z |= 4'b0100; 
	if(x==?20'b??1?1?00?011??001?01) z |= 4'b1000; 
	if(x==?20'b?1??1?00?011??001?01) z |= 4'b1000; 
	if(x==?20'b11????10?101?010?10?) z |= 4'b1000; 
	if(x==?20'b11????1?1101?101?10?) z |= 4'b1000; 
	if(x==?20'b1????10???00?1110?11) z |= 4'b1000; 
	if(x==?20'b??11?1??1011101??10?) z |= 4'b0100; 
	if(x==?20'b??1?1?001?0??1101?11) z |= 4'b1000; 
	if(x==?20'b1???1?001110?0?01??1) z |= 4'b1000; 
	if(x==?20'b?1??001?111??00?0?01) z |= 4'b0100; 
	if(x==?20'b?1??00?1?0?1011?1?11) z |= 4'b0100; 
	if(x==?20'b???100?101110?0?1??1) z |= 4'b0100; 
	if(x==?20'b??1??100?111?00?0?01) z |= 4'b1000; 
	if(x==?20'b?11?00??1011?1??011?) z |= 4'b0100; 
	if(x==?20'b??111???010?010?110?) z |= 4'b0100; 
	if(x==?20'b????0111?111110?10??) z |= 4'b0100; 
	if(x==?20'b?11???001101??1?011?) z |= 4'b1000; 
	if(x==?20'b?1???01?111?000?0?01) z |= 4'b0100; 
	if(x==?20'b111????1??01?0?11100) z |= 4'b1000; 
	if(x==?20'b111????1?0?1??011100) z |= 4'b1000; 
	if(x==?20'b????1110111??01110??) z |= 4'b1000; 
	if(x==?20'b??1??10??111?0000?01) z |= 4'b1000; 
	if(x==?20'b1?1?1?111110?0?01?1?) z |= 4'b1000; 
	if(x==?20'b?1??1?11100??11?1?01) z |= 4'b1000; 
	if(x==?20'b????1011010??1??010?) z |= 4'b0100; 
	if(x==?20'b?1?10??1111??00?0?01) z |= 4'b0100; 
	if(x==?20'b?1?111?101110?0?1?1?) z |= 4'b0100; 
	if(x==?20'b11?????1?010?010110?) z |= 4'b1000; 
	if(x==?20'b1?1?1??0?111?00?0?01) z |= 4'b1000; 
	if(x==?20'b??1?11?1?001?11?1?01) z |= 4'b0100; 
	if(x==?20'b?1?111?111?1?00?1?10) z |= 4'b0100; 
	if(x==?20'b1?1?1?111?11?00?1?10) z |= 4'b1000; 
	if(x==?20'b?1?1???1111?000?0?01) z |= 4'b0100; 
	if(x==?20'b?1?1?01?111??00?0?01) z |= 4'b0100; 
	if(x==?20'b??1?1?0?1110?1101?1?) z |= 4'b1000; 
	if(x==?20'b?1??1?0?1110?1101?1?) z |= 4'b1000; 
	if(x==?20'b1?1?1????111?0000?01) z |= 4'b1000; 
	if(x==?20'b?11???10?101?101?10?) z |= 4'b1000; 
	if(x==?20'b?11?01??101?101??10?) z |= 4'b0100; 
	if(x==?20'b??1??0?10111011?1?1?) z |= 4'b0100; 
	if(x==?20'b?1???0?10111011?1?1?) z |= 4'b0100; 
	if(x==?20'b1?1??10??111?00?0?01) z |= 4'b1000; 
	if(x==?20'b?1??00?1?0?1110?1?11) z |= 4'b0100; 
	if(x==?20'b??1?1?001?0??0111?11) z |= 4'b1000; 
	if(x==?20'b???10?1?0111011?1?1?) z |= 4'b0100; 
	if(x==?20'b??11?1??1011010??10?) z |= 4'b0100; 
	if(x==?20'b11????1?1101?010?10?) z |= 4'b1000; 
	if(x==?20'b?1111???10???10?1100) z |= 4'b0100; 
	if(x==?20'b???10?1?110100??1?01) z |= 4'b0100; 
	if(x==?20'b???100?1010??1???110) z |= 4'b0100; 
	if(x==?20'b1????1?01011??001?01) z |= 4'b1000; 
	if(x==?20'b111???1??101?101?10?) z |= 4'b1000; 
	if(x==?20'b?111?1??101?101??10?) z |= 4'b0100; 
	if(x==?20'b11?????01101?101?11?) z |= 4'b1000; 
	if(x==?20'b?1110???010?101??11?) z |= 4'b0100; 
	if(x==?20'b??1?00?1110??00?1?01) z |= 4'b0100; 
	if(x==?20'b1???1?00?010??1??110) z |= 4'b1000; 
	if(x==?20'b?1??00?1110??00?1?01) z |= 4'b0100; 
	if(x==?20'b??110???1011101??11?) z |= 4'b0100; 
	if(x==?20'b??1??0?10111110?1?1?) z |= 4'b0100; 
	if(x==?20'b?1???0?10111110?1?1?) z |= 4'b0100; 
	if(x==?20'b111????0?010?101?11?) z |= 4'b1000; 
	if(x==?20'b??1?1?00?011?00?1?01) z |= 4'b1000; 
	if(x==?20'b?1??1?00?011?00?1?01) z |= 4'b1000; 
	if(x==?20'b??1?1?0?1110?0111?1?) z |= 4'b1000; 
	if(x==?20'b?1??1?0?1110?0111?1?) z |= 4'b1000; 
	if(x==?20'b??1??0?1110?000?1?01) z |= 4'b0100; 
	if(x==?20'b?1???0?1110?000?1?01) z |= 4'b0100; 
	if(x==?20'b???1111?00??111???01) z |= 4'b0100; 
	if(x==?20'b1?1?1??01?0??1101?11) z |= 4'b1000; 
	if(x==?20'b???10?1?0111110?1?1?) z |= 4'b0100; 
	if(x==?20'b??1?1?0??011?0001?01) z |= 4'b1000; 
	if(x==?20'b?1??1?0??011?0001?01) z |= 4'b1000; 
	if(x==?20'b?1??1??01110?1101?1?) z |= 4'b1000; 
	if(x==?20'b????1011101?1?1?01??) z |= 4'b0100; 
	if(x==?20'b1????111??00?111??01) z |= 4'b1000; 
	if(x==?20'b????1101?101?1?101??) z |= 4'b1000; 
	if(x==?20'b?1?10??1?0?1011?1?11) z |= 4'b0100; 
	if(x==?20'b??1?0??10111011?1?1?) z |= 4'b0100; 
	if(x==?20'b??1?1?00??11?0001?01) z |= 4'b1000; 
	if(x==?20'b?11?01??101?010??10?) z |= 4'b0100; 
	if(x==?20'b?1???01?00??111?0?11) z |= 4'b0100; 
	if(x==?20'b?11111?1011?0?0?1?1?) z |= 4'b0100; 
	if(x==?20'b111?1?11?110?0?01?1?) z |= 4'b1000; 
	if(x==?20'b?1111???100??01?11?0) z |= 4'b0100; 
	if(x==?20'b????11?1?010??10010?) z |= 4'b1000; 
	if(x==?20'b??1?001??0??111?0?11) z |= 4'b0100; 
	if(x==?20'b?11???10?101?010?10?) z |= 4'b1000; 
	if(x==?20'b111???111110?0?01?1?) z |= 4'b1000; 
	if(x==?20'b?11???1?1101?101?10?) z |= 4'b1000; 
	if(x==?20'b??1??10???00?1110?11) z |= 4'b1000; 
	if(x==?20'b?11101??0111?1???10?) z |= 4'b0100; 
	if(x==?20'b1???1??01?00?111??11) z |= 4'b1000; 
	if(x==?20'b???10??100?1111???11) z |= 4'b0100; 
	if(x==?20'b?11111??01110?0?1?1?) z |= 4'b0100; 
	if(x==?20'b??1?0??1110100??1?01) z |= 4'b0100; 
	if(x==?20'b?1???100??0??1110?11) z |= 4'b1000; 
	if(x==?20'b111???101110??1??10?) z |= 4'b1000; 
	if(x==?20'b?11??1??1011101??10?) z |= 4'b0100; 
	if(x==?20'b?1??1??01011??001?01) z |= 4'b1000; 
	if(x==?20'b?11?01100000?0??1?1?) z |= 4'b1100; 
	if(x==?20'b?11?01100000??0?1?1?) z |= 4'b1100; 
	if(x==?20'b?1?1???100??111?0?11) z |= 4'b0100; 
	if(x==?20'b??1?1?001110?0?01??1) z |= 4'b1000; 
	if(x==?20'b???111??000?11??1?01) z |= 4'b0100; 
	if(x==?20'b1?1?1?????00?1110?11) z |= 4'b1000; 
	if(x==?20'b?1??00?101110?0?1??1) z |= 4'b0100; 
	if(x==?20'b111???11??00?1101??1) z |= 4'b1000; 
	if(x==?20'b????111?00?1111???01) z |= 4'b0100; 
	if(x==?20'b?11?1???010?010?110?) z |= 4'b0100; 
	if(x==?20'b?????1111?00?111??01) z |= 4'b1000; 
	if(x==?20'b??1???110000?11?1?01) z |= 4'b1100; 
	if(x==?20'b?1????110000?11?1?01) z |= 4'b1100; 
	if(x==?20'b?1?10??1?0?1110?1?11) z |= 4'b0100; 
	if(x==?20'b?11111?11101?0??1?1?) z |= 4'b0100; 
	if(x==?20'b1?????11?000??111?01) z |= 4'b1000; 
	if(x==?20'b?1110???010?010??11?) z |= 4'b0100; 
	if(x==?20'b??1?0??10111110?1?1?) z |= 4'b0100; 
	if(x==?20'b111?1?111011??0?1?1?) z |= 4'b1000; 
	if(x==?20'b??110???1011010??11?) z |= 4'b0100; 
	if(x==?20'b1?1?1??01?0??0111?11) z |= 4'b1000; 
	if(x==?20'b11?????01101?010?11?) z |= 4'b1000; 
	if(x==?20'b????0?1?1101000?1?01) z |= 4'b0100; 
	if(x==?20'b?11????1?010?010110?) z |= 4'b1000; 
	if(x==?20'b??110???100?010?111?) z |= 4'b0100; 
	if(x==?20'b?1??1??01110?0111?1?) z |= 4'b1000; 
	if(x==?20'b?11101??011??10??10?) z |= 4'b0100; 
	if(x==?20'b????1?1101??101?010?) z |= 4'b0100; 
	if(x==?20'b?????1?01011?0001?01) z |= 4'b1000; 
	if(x==?20'b111????0?010?010?11?) z |= 4'b1000; 
	if(x==?20'b?????11?010?101?010?) z |= 4'b0100; 
	if(x==?20'b1?1????0?001?100111?) z |= 4'b1000; 
	if(x==?20'b?1?10???100?001?111?) z |= 4'b0100; 
	if(x==?20'b111???10?110?01??10?) z |= 4'b1000; 
	if(x==?20'b?1110???101?101??11?) z |= 4'b0100; 
	if(x==?20'b111????0?101?101?11?) z |= 4'b1000; 
	if(x==?20'b?????11??010?101010?) z |= 4'b1000; 
	if(x==?20'b111????01?10?101?11?) z |= 4'b1000; 
	if(x==?20'b?1110???01?1101??11?) z |= 4'b0100; 
	if(x==?20'b?111?1??011?010??10?) z |= 4'b0100; 
	if(x==?20'b11?????0?001?010111?) z |= 4'b1000; 
	if(x==?20'b????0111010??1??010?) z |= 4'b0100; 
	if(x==?20'b111???1??110?010?10?) z |= 4'b1000; 
	if(x==?20'b????11??000111??1?01) z |= 4'b0100; 
	if(x==?20'b???10?1?1101?00?1?01) z |= 4'b0100; 
	if(x==?20'b???1?1??000?101??101) z |= 4'b0100; 
	if(x==?20'b1?????1??000?101?101) z |= 4'b1000; 
	if(x==?20'b1?1??1?01??0?1101?11) z |= 4'b1000; 
	if(x==?20'b?????111010?01??010?) z |= 4'b0100; 
	if(x==?20'b????1110?010??1?010?) z |= 4'b1000; 
	if(x==?20'b?1?10?1?0??1011?1?11) z |= 4'b0100; 
	if(x==?20'b1????1?01011?00?1?01) z |= 4'b1000; 
	if(x==?20'b?1??0?1?0111011?1?1?) z |= 4'b0100; 
	if(x==?20'b????0111?10?01??010?) z |= 4'b0100; 
	if(x==?20'b??????111000??111?01) z |= 4'b1000; 
	if(x==?20'b?11??1??1011010??10?) z |= 4'b0100; 
	if(x==?20'b???1??1?1101000?1?01) z |= 4'b0100; 
	if(x==?20'b?11???1?1101?010?10?) z |= 4'b1000; 
	if(x==?20'b??110???010?001?111?) z |= 4'b0100; 
	if(x==?20'b11?????0?010?100111?) z |= 4'b1000; 
	if(x==?20'b?1110???101101???11?) z |= 4'b0100; 
	if(x==?20'b1????1??1011?0001?01) z |= 4'b1000; 
	if(x==?20'b111???11??00?0111??1) z |= 4'b1000; 
	if(x==?20'b????1110?01???10010?) z |= 4'b1000; 
	if(x==?20'b111????01101??10?11?) z |= 4'b1000; 
	if(x==?20'b???111??000??11?1?01) z |= 4'b0100; 
	if(x==?20'b?1??0?1?110100??1?01) z |= 4'b0100; 
	if(x==?20'b??1?0?1?11010?0?1?01) z |= 4'b0100; 
	if(x==?20'b?1??00?1010??1???110) z |= 4'b0100; 
	if(x==?20'b1?????11?000?11?1?01) z |= 4'b1000; 
	if(x==?20'b?1?10??111??000?1?01) z |= 4'b0100; 
	if(x==?20'b?1???1?01011?0?01?01) z |= 4'b1000; 
	if(x==?20'b????101?011101??01??) z |= 4'b0100; 
	if(x==?20'b??1??1?01011??001?01) z |= 4'b1000; 
	if(x==?20'b?1?10???100?100?111?) z |= 4'b0100; 
	if(x==?20'b1?1?1??0??11?0001?01) z |= 4'b1000; 
	if(x==?20'b?11????01101?101?11?) z |= 4'b1000; 
	if(x==?20'b?1110???100?0?1?111?) z |= 4'b0100; 
	if(x==?20'b???111?100??11??1?01) z |= 4'b0100; 
	if(x==?20'b???100?1011?11??1?1?) z |= 4'b0100; 
	if(x==?20'b?????1011110??1001??) z |= 4'b1000; 
	if(x==?20'b11?????01?00?111??11) z |= 4'b1000; 
	if(x==?20'b??1?1?00?010??1??110) z |= 4'b1000; 
	if(x==?20'b?11?0???1011101??11?) z |= 4'b0100; 
	if(x==?20'b111?1?11??0??1101??1) z |= 4'b1000; 
	if(x==?20'b111????0?001??10111?) z |= 4'b1000; 
	if(x==?20'b?11111?1?0??011?1??1) z |= 4'b0100; 
	if(x==?20'b1?1????0?001?001111?) z |= 4'b1000; 
	if(x==?20'b1?1??1??1110?1101?1?) z |= 4'b1000; 
	if(x==?20'b111???111?0??1101??1) z |= 4'b1000; 
	if(x==?20'b??????1?1000?101?101) z |= 4'b1000; 
	if(x==?20'b?1?1??1?0111011?1?1?) z |= 4'b0100; 
	if(x==?20'b?1?10?1?1101?0??1?01) z |= 4'b0100; 
	if(x==?20'b????11?1?010?01?010?) z |= 4'b1000; 
	if(x==?20'b1???1?11??00??111?01) z |= 4'b1000; 
	if(x==?20'b?????1??0001101??101) z |= 4'b0100; 
	if(x==?20'b?1??111?00??111???01) z |= 4'b0100; 
	if(x==?20'b?1?10?1?0??1110?1?11) z |= 4'b0100; 
	if(x==?20'b?11111???0?1011?1??1) z |= 4'b0100; 
	if(x==?20'b1?1??1?01011??0?1?01) z |= 4'b1000; 
	if(x==?20'b??1?0??11101?00?1?01) z |= 4'b0100; 
	if(x==?20'b?1??0?1?0111110?1?1?) z |= 4'b0100; 
	if(x==?20'b?????11?010?010?010?) z |= 4'b0100; 
	if(x==?20'b1?1?1??01110?0?01??1) z |= 4'b1000; 
	if(x==?20'b?1??1??01011?00?1?01) z |= 4'b1000; 
	if(x==?20'b?11100?111??0?0?1??1) z |= 4'b0100; 
	if(x==?20'b??110???010?100?111?) z |= 4'b0100; 
	if(x==?20'b??1??111??00?111??01) z |= 4'b1000; 
	if(x==?20'b?1?1??1?110100??1?01) z |= 4'b0100; 
	if(x==?20'b?1110???101?010??11?) z |= 4'b0100; 
	if(x==?20'b1?1??1?01??0?0111?11) z |= 4'b1000; 
	if(x==?20'b?1?10??101110?0?1??1) z |= 4'b0100; 
	if(x==?20'b?1110???01?1010??11?) z |= 4'b0100; 
	if(x==?20'b111?1?00??11?0?01??1) z |= 4'b1000; 
	if(x==?20'b???1111?111?000???10) z |= 4'b0100; 
	if(x==?20'b1?1??1??1011??001?01) z |= 4'b1000; 
	if(x==?20'b????11?1??10?010010?) z |= 4'b1000; 
	if(x==?20'b??1????11101000?1?01) z |= 4'b0100; 
	if(x==?20'b?????111?10?101?010?) z |= 4'b0100; 
	if(x==?20'b?111011?11??011?1???) z |= 4'b0100; 
	if(x==?20'b??????111000?11?1?01) z |= 4'b1000; 
	if(x==?20'b111????0?101?010?11?) z |= 4'b1000; 
	if(x==?20'b????111??01??101010?) z |= 4'b1000; 
	if(x==?20'b?1??1???1011?0001?01) z |= 4'b1000; 
	if(x==?20'b111?????1101?101?11?) z |= 4'b1000; 
	if(x==?20'b?????11??010?010010?) z |= 4'b1000; 
	if(x==?20'b111????01?10?010?11?) z |= 4'b1000; 
	if(x==?20'b1????111?111?000??10) z |= 4'b1000; 
	if(x==?20'b????11??0001?11?1?01) z |= 4'b0100; 
	if(x==?20'b11?????0?010?001111?) z |= 4'b1000; 
	if(x==?20'b???1?1??000?010??101) z |= 4'b0100; 
	if(x==?20'b??1?1??01?00?111??11) z |= 4'b1000; 
	if(x==?20'b?111????1011101??11?) z |= 4'b0100; 
	if(x==?20'b?1??0??100?1111???11) z |= 4'b0100; 
	if(x==?20'b111??110??11?1101???) z |= 4'b1000; 
	if(x==?20'b?11111??0?1?011?1??1) z |= 4'b0100; 
	if(x==?20'b1?????1??000?010?101) z |= 4'b1000; 
	if(x==?20'b????1011?11?101?01??) z |= 4'b0100; 
	if(x==?20'b????1101?11??10101??) z |= 4'b1000; 
	if(x==?20'b?11111?1?0??110?1??1) z |= 4'b0100; 
	if(x==?20'b??1?11??000?11??1?01) z |= 4'b0100; 
	if(x==?20'b?1??11??000?11??1?01) z |= 4'b0100; 
	if(x==?20'b111????0?001?0?1111?) z |= 4'b1000; 
	if(x==?20'b??1?11?11101?00?1?10) z |= 4'b1100; 
	if(x==?20'b?1?1??1?0111110?1?1?) z |= 4'b0100; 
	if(x==?20'b??11111??0??111???01) z |= 4'b0100; 
	if(x==?20'b?1??1?111011?00?1?10) z |= 4'b1100; 
	if(x==?20'b?11111???0?1110?1??1) z |= 4'b0100; 
	if(x==?20'b1?1?????1100?010111?) z |= 4'b1000; 
	if(x==?20'b?1?1????0011010?111?) z |= 4'b0100; 
	if(x==?20'b111?1?11??0??0111??1) z |= 4'b1000; 
	if(x==?20'b11???111??0??111??01) z |= 4'b1000; 
	if(x==?20'b????1?001?00?11?1?11) z |= 4'b1000; 
	if(x==?20'b1?1??1??1110?0111?1?) z |= 4'b1000; 
	if(x==?20'b???10?110??1111???11) z |= 4'b0100; 
	if(x==?20'b111???111?0??0111??1) z |= 4'b1000; 
	if(x==?20'b???10??1010?00???101) z |= 4'b0100; 
	if(x==?20'b1???1?11??00?11?1?01) z |= 4'b1000; 
	if(x==?20'b1???11?01??0?111??11) z |= 4'b1000; 
	if(x==?20'b???111?100???11?1?01) z |= 4'b0100; 
	if(x==?20'b??1???11?000??111?01) z |= 4'b1000; 
	if(x==?20'b?1????11?000??111?01) z |= 4'b1000; 
	if(x==?20'b1???1?00?110?11?1?1?) z |= 4'b1000; 
	if(x==?20'b????00?100?1?11?1?11) z |= 4'b0100; 
	if(x==?20'b?11?0???1011010??11?) z |= 4'b0100; 
	if(x==?20'b?1?1111?111?00????10) z |= 4'b0100; 
	if(x==?20'b1???1??0?010??00?101) z |= 4'b1000; 
	if(x==?20'b??11111?111?0?0???10) z |= 4'b0100; 
	if(x==?20'b?11????01101?010?11?) z |= 4'b1000; 
	if(x==?20'b?111011?11??110?1???) z |= 4'b0100; 
	if(x==?20'b????1?0?1?00?1101?11) z |= 4'b1000; 
	if(x==?20'b11??1??01?0??111??11) z |= 4'b1000; 
	if(x==?20'b?11?0???100?010?111?) z |= 4'b0100; 
	if(x==?20'b11???111?111?0?0??10) z |= 4'b1000; 
	if(x==?20'b1?1??111?111??00??10) z |= 4'b1000; 
	if(x==?20'b?????111010??10?010?) z |= 4'b0100; 
	if(x==?20'b?????0?100?1011?1?11) z |= 4'b0100; 
	if(x==?20'b?11111??0?1?110?1??1) z |= 4'b0100; 
	if(x==?20'b?1??11?01?11?0111?1?) z |= 4'b1000; 
	if(x==?20'b?????1??0001010??101) z |= 4'b0100; 
	if(x==?20'b??????1?1000?010?101) z |= 4'b1000; 
	if(x==?20'b?????1?11101?10101??) z |= 4'b1000; 
	if(x==?20'b???100?1?11?011?1?1?) z |= 4'b0100; 
	if(x==?20'b????0111?10??10?010?) z |= 4'b0100; 
	if(x==?20'b????1?1?1011101?01??) z |= 4'b0100; 
	if(x==?20'b????011101???10?010?) z |= 4'b0100; 
	if(x==?20'b?11????0?001?010111?) z |= 4'b1000; 
	if(x==?20'b?????1101?10?10101??) z |= 4'b1000; 
	if(x==?20'b????011?01?1101?01??) z |= 4'b0100; 
	if(x==?20'b111??110??11?0111???) z |= 4'b1000; 
	if(x==?20'b?1110???1011?10??11?) z |= 4'b0100; 
	if(x==?20'b????1110?01??01?010?) z |= 4'b1000; 
	if(x==?20'b111????01101?01??11?) z |= 4'b1000; 
	if(x==?20'b?111??1?011?011?1?1?) z |= 4'b0100; 
	if(x==?20'b????1101?1?1?01001??) z |= 4'b1000; 
	if(x==?20'b????1110??10?01?010?) z |= 4'b1000; 
	if(x==?20'b1???1?0?1?00?11?1?11) z |= 4'b1000; 
	if(x==?20'b?1??0?1?1101?00?1?01) z |= 4'b0100; 
	if(x==?20'b?????111?10?010?010?) z |= 4'b0100; 
	if(x==?20'b111??1???110?1101?1?) z |= 4'b1000; 
	if(x==?20'b?1???1??000?101??101) z |= 4'b0100; 
	if(x==?20'b1???1??0??00?1101?11) z |= 4'b1000; 
	if(x==?20'b??1???1??000?101?101) z |= 4'b1000; 
	if(x==?20'b??1?111??0?1111???01) z |= 4'b0100; 
	if(x==?20'b???10??100??011?1?11) z |= 4'b0100; 
	if(x==?20'b?1110???100??10?111?) z |= 4'b0100; 
	if(x==?20'b1?????101?00?101?1?1) z |= 4'b1000; 
	if(x==?20'b?1???1111?0??111??01) z |= 4'b1000; 
	if(x==?20'b??1??1?01011?00?1?01) z |= 4'b1000; 
	if(x==?20'b????101?0111?10?01??) z |= 4'b0100; 
	if(x==?20'b???1?0?100?1?11?1?11) z |= 4'b0100; 
	if(x==?20'b1??????01?00?1101?11) z |= 4'b1000; 
	if(x==?20'b?111????1011010??11?) z |= 4'b0100; 
	if(x==?20'b????111??01??010010?) z |= 4'b1000; 
	if(x==?20'b???101??00?1101??1?1) z |= 4'b0100; 
	if(x==?20'b111?????1101?010?11?) z |= 4'b1000; 
	if(x==?20'b?1????1?1101000?1?01) z |= 4'b0100; 
	if(x==?20'b???10???00?1011?1?11) z |= 4'b0100; 
	if(x==?20'b?????1011110?01?01??) z |= 4'b1000; 
	if(x==?20'b?11?0???010?001?111?) z |= 4'b0100; 
	if(x==?20'b?11????0?010?100111?) z |= 4'b1000; 
	if(x==?20'b??110???0?11111???11) z |= 4'b0100; 
	if(x==?20'b????1011?11?010?01??) z |= 4'b0100; 
	if(x==?20'b??1??1??1011?0001?01) z |= 4'b1000; 
	if(x==?20'b??1?11??000??11?1?01) z |= 4'b0100; 
	if(x==?20'b?1??11??000??11?1?01) z |= 4'b0100; 
	if(x==?20'b????0111011??11?10??) z |= 4'b0100; 
	if(x==?20'b????1110?110?11?10??) z |= 4'b1000; 
	if(x==?20'b?1?10??111?1000?1??1) z |= 4'b0100; 
	if(x==?20'b?????0?100?1110?1?11) z |= 4'b0100; 
	if(x==?20'b1?1?1??01?11?0001??1) z |= 4'b1000; 
	if(x==?20'b??1?0??1111?00??0?01) z |= 4'b0100; 
	if(x==?20'b??1?001?111??0??0?01) z |= 4'b0100; 
	if(x==?20'b????1?0?1?00?0111?11) z |= 4'b1000; 
	if(x==?20'b??1?11?100??11??1?01) z |= 4'b0100; 
	if(x==?20'b?1??11?100??11??1?01) z |= 4'b0100; 
	if(x==?20'b?1??1??0?111??000?01) z |= 4'b1000; 
	if(x==?20'b?11????01?00?111??11) z |= 4'b1000; 
	if(x==?20'b?1?1??1?1101?00?1?01) z |= 4'b0100; 
	if(x==?20'b?????111011?011?10??) z |= 4'b0100; 
	if(x==?20'b????111??110?11010??) z |= 4'b1000; 
	if(x==?20'b??1?11?111?100??1?10) z |= 4'b0100; 
	if(x==?20'b????0111011?01??01??) z |= 4'b0100; 
	if(x==?20'b?1??1?111?11??001?10) z |= 4'b1000; 
	if(x==?20'b?1???100?111??0?0?01) z |= 4'b1000; 
	if(x==?20'b1?1??1??1011?00?1?01) z |= 4'b1000; 
	if(x==?20'b?111??1?011?110?1?1?) z |= 4'b0100; 
	if(x==?20'b1???1?00?11??0111?1?) z |= 4'b1000; 
	if(x==?20'b????1??01?00?1101?11) z |= 4'b1000; 
	if(x==?20'b?1?11???100?000?111?) z |= 4'b0100; 
	if(x==?20'b????1110?110??1001??) z |= 4'b1000; 
	if(x==?20'b??1??01?111?00??0?01) z |= 4'b0100; 
	if(x==?20'b???10??100??110?1?11) z |= 4'b0100; 
	if(x==?20'b??1?1?11??00??111?01) z |= 4'b1000; 
	if(x==?20'b?1??1?11??00??111?01) z |= 4'b1000; 
	if(x==?20'b??1?1?00?110??111?1?) z |= 4'b1000; 
	if(x==?20'b????0??100?1011?1?11) z |= 4'b0100; 
	if(x==?20'b1?1????1?001?000111?) z |= 4'b1000; 
	if(x==?20'b?1???10??111??000?01) z |= 4'b1000; 
	if(x==?20'b?1?10?110???111???11) z |= 4'b0100; 
	if(x==?20'b111????0?01??100111?) z |= 4'b1000; 
	if(x==?20'b111????0??10?100111?) z |= 4'b1000; 
	if(x==?20'b?1110????10?001?111?) z |= 4'b0100; 
	if(x==?20'b???10???00?1110?1?11) z |= 4'b0100; 
	if(x==?20'b????0??1010?000??101) z |= 4'b0100; 
	if(x==?20'b?11?0???010?100?111?) z |= 4'b0100; 
	if(x==?20'b111??1???110?0111?1?) z |= 4'b1000; 
	if(x==?20'b????1?1?1011010?01??) z |= 4'b0100; 
	if(x==?20'b1???1??0??00?0111?11) z |= 4'b1000; 
	if(x==?20'b?1110???0?1?001?111?) z |= 4'b0100; 
	if(x==?20'b1?1?11?0???0?111??11) z |= 4'b1000; 
	if(x==?20'b????1??0?010?000?101) z |= 4'b1000; 
	if(x==?20'b??110?1?0??1111???11) z |= 4'b0100; 
	if(x==?20'b?1??111?111?000???10) z |= 4'b0100; 
	if(x==?20'b?1?10?1??0?1111???11) z |= 4'b0100; 
	if(x==?20'b????011?01?1010?01??) z |= 4'b0100; 
	if(x==?20'b1?1??1?01?0??111??11) z |= 4'b1000; 
	if(x==?20'b?????1?11101?01001??) z |= 4'b1000; 
	if(x==?20'b1??????01?00?0111?11) z |= 4'b1000; 
	if(x==?20'b11???1?01??0?111??11) z |= 4'b1000; 
	if(x==?20'b111??1??1110?11?1?1?) z |= 4'b1000; 
	if(x==?20'b????11101?1??10101??) z |= 4'b1000; 
	if(x==?20'b??1??111?111?000??10) z |= 4'b1000; 
	if(x==?20'b?111??1?0111?11?1?1?) z |= 4'b0100; 
	if(x==?20'b?????1101?10?01001??) z |= 4'b1000; 
	if(x==?20'b?11????0?010?001111?) z |= 4'b1000; 
	if(x==?20'b?1???1??000?010??101) z |= 4'b0100; 
	if(x==?20'b??111???010?000?111?) z |= 4'b0100; 
	if(x==?20'b?1110??111?10?0?1??1) z |= 4'b0100; 
	if(x==?20'b111?1??01?11?0?01??1) z |= 4'b1000; 
	if(x==?20'b????0111?1?1101?01??) z |= 4'b0100; 
	if(x==?20'b???100?1011?00??1??1) z |= 4'b0100; 
	if(x==?20'b??1???1??000?010?101) z |= 4'b1000; 
	if(x==?20'b1???1?00?110??001??1) z |= 4'b1000; 
	if(x==?20'b???101??00?1010??1?1) z |= 4'b0100; 
	if(x==?20'b??1101??1011?1???10?) z |= 4'b0100; 
	if(x==?20'b1???1???1?00?1101?11) z |= 4'b1000; 
	if(x==?20'b?????111011?110?10??) z |= 4'b0100; 
	if(x==?20'b11?????1?010?000111?) z |= 4'b1000; 
	if(x==?20'b???10??1010??00??101) z |= 4'b0100; 
	if(x==?20'b1?????101?00?010?1?1) z |= 4'b1000; 
	if(x==?20'b11????101101??1??10?) z |= 4'b1000; 
	if(x==?20'b1???1??0?010?00??101) z |= 4'b1000; 
	if(x==?20'b111????0?0?1?001111?) z |= 4'b1000; 
	if(x==?20'b?1?1111?111??00???10) z |= 4'b0100; 
	if(x==?20'b???1???100?1011?1?11) z |= 4'b0100; 
	if(x==?20'b?11?111??0??111???01) z |= 4'b0100; 
	if(x==?20'b?1111???100?0?0?111?) z |= 4'b0100; 
	if(x==?20'b1???1?111??0?0001?11) z |= 4'b1000; 
	if(x==?20'b????111??110?10101??) z |= 4'b1000; 
	if(x==?20'b1?1??111?111?00???10) z |= 4'b1000; 
	if(x==?20'b???1???1010?000??101) z |= 4'b0100; 
	if(x==?20'b??111???010?10??110?) z |= 4'b0100; 
	if(x==?20'b????111??110?01110??) z |= 4'b1000; 
	if(x==?20'b??110??1??11111???11) z |= 4'b0100; 
	if(x==?20'b????1?1??001?100110?) z |= 4'b1000; 
	if(x==?20'b????0??100?1110?1?11) z |= 4'b0100; 
	if(x==?20'b???111?10??1000?1?11) z |= 4'b0100; 
	if(x==?20'b111????1?001?0?0111?) z |= 4'b1000; 
	if(x==?20'b1???1????010?000?101) z |= 4'b1000; 
	if(x==?20'b?11??111??0??111??01) z |= 4'b1000; 
	if(x==?20'b???10??1?10?000??101) z |= 4'b0100; 
	if(x==?20'b?????1?1100?001?110?) z |= 4'b0100; 
	if(x==?20'b?1110????10?100?111?) z |= 4'b0100; 
	if(x==?20'b?1??0?110??1111???11) z |= 4'b0100; 
	if(x==?20'b????1??01?00?0111?11) z |= 4'b1000; 
	if(x==?20'b1???1??0?01??000?101) z |= 4'b1000; 
	if(x==?20'b????111?1110?11?10??) z |= 4'b1000; 
	if(x==?20'b?1??0??1010?00???101) z |= 4'b0100; 
	if(x==?20'b??1?1?11??00?11?1?01) z |= 4'b1000; 
	if(x==?20'b??1?11?01??0?111??11) z |= 4'b1000; 
	if(x==?20'b?1??1?11??00?11?1?01) z |= 4'b1000; 
	if(x==?20'b??1?11?100???11?1?01) z |= 4'b0100; 
	if(x==?20'b?1??11?100???11?1?01) z |= 4'b0100; 
	if(x==?20'b?1110???0?1?100?111?) z |= 4'b0100; 
	if(x==?20'b??1?00?1011??11?1?1?) z |= 4'b0100; 
	if(x==?20'b1???1100110????01?1?) z |= 4'b1000; 
	if(x==?20'b?1??00?1011??11?1?1?) z |= 4'b0100; 
	if(x==?20'b?1??1?00?110?11?1?1?) z |= 4'b1000; 
	if(x==?20'b?11?1???0100?01?110?) z |= 4'b1100; 
	if(x==?20'b?????1110111?11?10??) z |= 4'b0100; 
	if(x==?20'b??1?1??0?010??00?101) z |= 4'b1000; 
	if(x==?20'b?11?111?111?0?0???10) z |= 4'b0100; 
	if(x==?20'b11?????1?010??01110?) z |= 4'b1000; 
	if(x==?20'b?11?1??01?0??111??11) z |= 4'b1000; 
	if(x==?20'b111????0??10?001111?) z |= 4'b1000; 
	if(x==?20'b???10011?0110???1?1?) z |= 4'b0100; 
	if(x==?20'b?11??111?111?0?0??10) z |= 4'b1000; 
	if(x==?20'b???1010??1??000??110) z |= 4'b0100; 
	if(x==?20'b?1?1011111?10???1?1?) z |= 4'b0100; 
	if(x==?20'b1????010??1??000?110) z |= 4'b1000; 
	if(x==?20'b1?1?11101?11???01?1?) z |= 4'b1000; 
	if(x==?20'b?1111???010?00??111?) z |= 4'b0100; 
	if(x==?20'b??1?1?00?11??1101?1?) z |= 4'b1000; 
	if(x==?20'b????1?001110??001??1) z |= 4'b1000; 
	if(x==?20'b????00?1011100??1??1) z |= 4'b0100; 
	if(x==?20'b1?1?1?0?100??0?011??) z |= 4'b1000; 
	if(x==?20'b111????1?010??00111?) z |= 4'b1000; 
	if(x==?20'b???10?11111?0?0???01) z |= 4'b0100; 
	if(x==?20'b???1???100?1110?1?11) z |= 4'b0100; 
	if(x==?20'b1???11?0?111?0?0??01) z |= 4'b1000; 
	if(x==?20'b1?1?1?111?0??0?01?11) z |= 4'b1000; 
	if(x==?20'b111?????1?10?100111?) z |= 4'b1000; 
	if(x==?20'b?1?1?0?1?0010?0?11??) z |= 4'b0100; 
	if(x==?20'b??1?1?0?1?00?11?1?11) z |= 4'b1000; 
	if(x==?20'b?1?1??110??1111???11) z |= 4'b0100; 
	if(x==?20'b??1?1??0??00?1101?11) z |= 4'b1000; 
	if(x==?20'b1???1???1?00?0111?11) z |= 4'b1000; 
	if(x==?20'b1?1?1?111??0??001?11) z |= 4'b1000; 
	if(x==?20'b?1??0??100??011?1?11) z |= 4'b0100; 
	if(x==?20'b1?1?11??1??0?111??11) z |= 4'b1000; 
	if(x==?20'b??1???101?00?101?1?1) z |= 4'b1000; 
	if(x==?20'b1???1???1101?101?11?) z |= 4'b1000; 
	if(x==?20'b?1??1?111110?0?01?1?) z |= 4'b1000; 
	if(x==?20'b?1?111?10??100??1?11) z |= 4'b0100; 
	if(x==?20'b?1???0?100?1?11?1?11) z |= 4'b0100; 
	if(x==?20'b?1?111?1?0?10?0?1?11) z |= 4'b0100; 
	if(x==?20'b??110?11???1111???11) z |= 4'b0100; 
	if(x==?20'b??1????01?00?1101?11) z |= 4'b1000; 
	if(x==?20'b?1?????01?00?1101?11) z |= 4'b1000; 
	if(x==?20'b11??11?01????111??11) z |= 4'b1000; 
	if(x==?20'b?????1?1100?100?110?) z |= 4'b0100; 
	if(x==?20'b????0111?1?1010?01??) z |= 4'b0100; 
	if(x==?20'b?111????0?11001?111?) z |= 4'b0100; 
	if(x==?20'b??1?0??1111??00?0?01) z |= 4'b0100; 
	if(x==?20'b??11???1010?101??11?) z |= 4'b0100; 
	if(x==?20'b?1??01??00?1101??1?1) z |= 4'b0100; 
	if(x==?20'b1???1?001110??0?1??1) z |= 4'b1000; 
	if(x==?20'b????11101?1??01001??) z |= 4'b1000; 
	if(x==?20'b???1???11011101??11?) z |= 4'b0100; 
	if(x==?20'b??1?11?101110?0?1?1?) z |= 4'b0100; 
	if(x==?20'b??1?0???00?1011?1?11) z |= 4'b0100; 
	if(x==?20'b?1??0???00?1011?1?11) z |= 4'b0100; 
	if(x==?20'b?1??1??0?111?00?0?01) z |= 4'b1000; 
	if(x==?20'b?11?0???0?11111???11) z |= 4'b0100; 
	if(x==?20'b11??1????010?101?11?) z |= 4'b1000; 
	if(x==?20'b???100?10111?0??1??1) z |= 4'b0100; 
	if(x==?20'b????1?1??001?001110?) z |= 4'b1000; 
	if(x==?20'b??1????1111?000?0?01) z |= 4'b0100; 
	if(x==?20'b1???1?0?1110??001??1) z |= 4'b1000; 
	if(x==?20'b??1??01?111??00?0?01) z |= 4'b0100; 
	if(x==?20'b?1??1????111?0000?01) z |= 4'b1000; 
	if(x==?20'b1?1?1??0??00?11?1?11) z |= 4'b1000; 
	if(x==?20'b???1?0?1011100??1??1) z |= 4'b0100; 
	if(x==?20'b??111???010??01?110?) z |= 4'b0100; 
	if(x==?20'b?????111011?010?01??) z |= 4'b0100; 
	if(x==?20'b?1?10??100???11?1?11) z |= 4'b0100; 
	if(x==?20'b?11111??110?00??1?1?) z |= 4'b0100; 
	if(x==?20'b11?????1?010?10?110?) z |= 4'b1000; 
	if(x==?20'b?1???10??111?00?0?01) z |= 4'b1000; 
	if(x==?20'b1?1?1?111110??0?1?1?) z |= 4'b1000; 
	if(x==?20'b??1?00?1?11?110?1?1?) z |= 4'b0100; 
	if(x==?20'b?1??00?1?11?110?1?1?) z |= 4'b0100; 
	if(x==?20'b????00?1011?000?1??1) z |= 4'b0100; 
	if(x==?20'b????1?00?110?0001??1) z |= 4'b1000; 
	if(x==?20'b1???1???1110?101?11?) z |= 4'b1000; 
	if(x==?20'b?1?111?10111?0??1?1?) z |= 4'b0100; 
	if(x==?20'b1????1?01?0??1101?11) z |= 4'b1000; 
	if(x==?20'b???1?1??010?000??110) z |= 4'b0100; 
	if(x==?20'b1?1?1?????00?1101?11) z |= 4'b1000; 
	if(x==?20'b???1???10111101??11?) z |= 4'b0100; 
	if(x==?20'b111???11?011??001?1?) z |= 4'b1000; 
	if(x==?20'b?1?10?11111?0?????01) z |= 4'b0100; 
	if(x==?20'b?1?1???100??011?1?11) z |= 4'b0100; 
	if(x==?20'b?????11?100?010?110?) z |= 4'b0100; 
	if(x==?20'b???10?1??0?1011?1?11) z |= 4'b0100; 
	if(x==?20'b1?????1??010?000?110) z |= 4'b1000; 
	if(x==?20'b?1??1?00?11??0111?1?) z |= 4'b1000; 
	if(x==?20'b???10?1?111?000???01) z |= 4'b0100; 
	if(x==?20'b1?1?11?0?111???0??01) z |= 4'b1000; 
	if(x==?20'b?1?1??1?0101010??1??) z |= 4'b0100; 
	if(x==?20'b?111?1??101?01???10?) z |= 4'b0100; 
	if(x==?20'b?111?1??01?101???10?) z |= 4'b0100; 
	if(x==?20'b?1??0??100??110?1?11) z |= 4'b0100; 
	if(x==?20'b?1?111?10???000?1?11) z |= 4'b0100; 
	if(x==?20'b??????101100?01011??) z |= 4'b1000; 
	if(x==?20'b1?1?1?11???0?0001?11) z |= 4'b1000; 
	if(x==?20'b1????1?0?111?000??01) z |= 4'b1000; 
	if(x==?20'b????01??0011010?11??) z |= 4'b0100; 
	if(x==?20'b1???1??01101?0?0?1?1) z |= 4'b1000; 
	if(x==?20'b?????11??001?010110?) z |= 4'b1000; 
	if(x==?20'b111???1??101??10?10?) z |= 4'b1000; 
	if(x==?20'b?111????0?11100?111?) z |= 4'b0100; 
	if(x==?20'b111???1?1?10??10?10?) z |= 4'b1000; 
	if(x==?20'b1?1??1??1010?010?1??) z |= 4'b1000; 
	if(x==?20'b111?????1?10?001111?) z |= 4'b1000; 
	if(x==?20'b???100?1011??00?1??1) z |= 4'b0100; 
	if(x==?20'b??1?0???00?1110?1?11) z |= 4'b0100; 
	if(x==?20'b?1??0???00?1110?1?11) z |= 4'b0100; 
	if(x==?20'b1???1?00?110?00?1??1) z |= 4'b1000; 
	if(x==?20'b???10??110110?0??1?1) z |= 4'b0100; 
	if(x==?20'b??1?1??0??00?0111?11) z |= 4'b1000; 
	if(x==?20'b?11111??011?00??1?1?) z |= 4'b0100; 
	if(x==?20'b?1?????11?01?100110?) z |= 4'b1000; 
	if(x==?20'b?11?0?1?0??1111???11) z |= 4'b0100; 
	if(x==?20'b111???11?110??001?1?) z |= 4'b1000; 
	if(x==?20'b??1????01?00?0111?11) z |= 4'b1000; 
	if(x==?20'b?1?????01?00?0111?11) z |= 4'b1000; 
	if(x==?20'b?11??1?01??0?111??11) z |= 4'b1000; 
	if(x==?20'b???1?0?1011?000?1??1) z |= 4'b0100; 
	if(x==?20'b1???1?0??110?0001??1) z |= 4'b1000; 
	if(x==?20'b?11?1???010?000?111?) z |= 4'b0100; 
	if(x==?20'b???100?1?11?000?1??1) z |= 4'b0100; 
	if(x==?20'b11???01?100???0011??) z |= 4'b1000; 
	if(x==?20'b?????1111111111???1?) z |= 4'b0100; 
	if(x==?20'b?1??00?1011?00??1??1) z |= 4'b0100; 
	if(x==?20'b??1?1?00?110??001??1) z |= 4'b1000; 
	if(x==?20'b??11???1010?010??11?) z |= 4'b0100; 
	if(x==?20'b?1??01??00?1010??1?1) z |= 4'b0100; 
	if(x==?20'b?11?01??1011?1???10?) z |= 4'b0100; 
	if(x==?20'b??1?1???1?00?1101?11) z |= 4'b1000; 
	if(x==?20'b?111101??1??101??1??) z |= 4'b0100; 
	if(x==?20'b?11????1?010?000111?) z |= 4'b1000; 
	if(x==?20'b????111?1111?111??1?) z |= 4'b1000; 
	if(x==?20'b?1??0??1010??00??101) z |= 4'b0100; 
	if(x==?20'b??1???101?00?010?1?1) z |= 4'b1000; 
	if(x==?20'b???1???11011010??11?) z |= 4'b0100; 
	if(x==?20'b1???1???1101?010?11?) z |= 4'b1000; 
	if(x==?20'b1???1100110??0??1?1?) z |= 4'b1000; 
	if(x==?20'b?11???101101??1??10?) z |= 4'b1000; 
	if(x==?20'b1???1100110???0?1?1?) z |= 4'b1000; 
	if(x==?20'b?1?1???100??110?1?11) z |= 4'b0100; 
	if(x==?20'b???10?1??0?1110?1?11) z |= 4'b0100; 
	if(x==?20'b?1??1??01?0??1101?11) z |= 4'b1000; 
	if(x==?20'b??1?1??0?010?00??101) z |= 4'b1000; 
	if(x==?20'b111??101??1??101?1??) z |= 4'b1000; 
	if(x==?20'b?1?????100?1011?1?11) z |= 4'b0100; 
	if(x==?20'b?1111???0?1?01??110?) z |= 4'b0100; 
	if(x==?20'b?1?10?1?111?00????01) z |= 4'b0100; 
	if(x==?20'b?????01?1110?10011??) z |= 4'b1000; 
	if(x==?20'b??110?1?111?0?0???01) z |= 4'b0100; 
	if(x==?20'b1???1??01110??001??1) z |= 4'b1000; 
	if(x==?20'b111????1?01??1?0110?) z |= 4'b1000; 
	if(x==?20'b11??1????010?010?11?) z |= 4'b1000; 
	if(x==?20'b??1?1?111??0?0001?11) z |= 4'b1000; 
	if(x==?20'b1????1?01?0??0111?11) z |= 4'b1000; 
	if(x==?20'b???10011?011?0??1?1?) z |= 4'b0100; 
	if(x==?20'b?1111????10?0?1?110?) z |= 4'b0100; 
	if(x==?20'b???10011?011??0?1?1?) z |= 4'b0100; 
	if(x==?20'b111????1??10?1?0110?) z |= 4'b1000; 
	if(x==?20'b???????01100?010111?) z |= 4'b1000; 
	if(x==?20'b?1?????1010?000??101) z |= 4'b0100; 
	if(x==?20'b?11?1???010?10??110?) z |= 4'b0100; 
	if(x==?20'b??1?0??1?0?1011?1?11) z |= 4'b0100; 
	if(x==?20'b????0???0011010?111?) z |= 4'b0100; 
	if(x==?20'b???10??1011100??1??1) z |= 4'b0100; 
	if(x==?20'b?11?0??1??11111???11) z |= 4'b0100; 
	if(x==?20'b1?1?11101?11?0??1?1?) z |= 4'b1000; 
	if(x==?20'b?1?1011111?1??0?1?1?) z |= 4'b0100; 
	if(x==?20'b1?1?1?????00?0111?11) z |= 4'b1000; 
	if(x==?20'b111????1?0?1?000111?) z |= 4'b1000; 
	if(x==?20'b?1??11?10??1000?1?11) z |= 4'b0100; 
	if(x==?20'b11???1?0?111?0?0??01) z |= 4'b1000; 
	if(x==?20'b?1111???010??00?111?) z |= 4'b0100; 
	if(x==?20'b1?1??1?0?111??00??01) z |= 4'b1000; 
	if(x==?20'b11??1????101?101?11?) z |= 4'b1000; 
	if(x==?20'b??1?1????010?000?101) z |= 4'b1000; 
	if(x==?20'b??11???1101?101??11?) z |= 4'b0100; 
	if(x==?20'b????1?001110?00?1??1) z |= 4'b1000; 
	if(x==?20'b?1??0??1?10?000??101) z |= 4'b0100; 
	if(x==?20'b11???11011???1101???) z |= 4'b1000; 
	if(x==?20'b111????111?0???1110?) z |= 4'b1000; 
	if(x==?20'b?????10?0111001?11??) z |= 4'b0100; 
	if(x==?20'b??1?1??0?01??000?101) z |= 4'b1000; 
	if(x==?20'b1??????01101?000?1?1) z |= 4'b1000; 
	if(x==?20'b????00?10111?00?1??1) z |= 4'b0100; 
	if(x==?20'b1?1?1???1?00?11?1?11) z |= 4'b1000; 
	if(x==?20'b111????1?010?00?111?) z |= 4'b1000; 
	if(x==?20'b??1?1100110????01?1?) z |= 4'b1000; 
	if(x==?20'b?1?1?11111?10?0?1?1?) z |= 4'b0100; 
	if(x==?20'b1?1?111?1?11?0?01?1?) z |= 4'b1000; 
	if(x==?20'b???10???1011000??1?1) z |= 4'b0100; 
	if(x==?20'b??11011???11011?1???) z |= 4'b0100; 
	if(x==?20'b???1???10111010??11?) z |= 4'b0100; 
	if(x==?20'b?11????1?010??01110?) z |= 4'b1000; 
	if(x==?20'b1???1???1110?010?11?) z |= 4'b1000; 
	if(x==?20'b?1?1???100?1?11?1?11) z |= 4'b0100; 
	if(x==?20'b????1?0?1110?0001??1) z |= 4'b1000; 
	if(x==?20'b?????100?001???1110?) z |= 4'b1001; 
	if(x==?20'b?1111????10?000?111?) z |= 4'b0100; 
	if(x==?20'b?1??0011?0110???1?1?) z |= 4'b0100; 
	if(x==?20'b1?1?1?111??0?00?1?11) z |= 4'b1000; 
	if(x==?20'b?????0?10111000?1??1) z |= 4'b0100; 
	if(x==?20'b?1111???01??000?111?) z |= 4'b0100; 
	if(x==?20'b?1??010??1??000??110) z |= 4'b0100; 
	if(x==?20'b??1??010??1??000?110) z |= 4'b1000; 
	if(x==?20'b?1?111?10??1?00?1?11) z |= 4'b0100; 
	if(x==?20'b??1????100??111?0?11) z |= 4'b0100; 
	if(x==?20'b?11111?1011??0??1?1?) z |= 4'b0100; 
	if(x==?20'b111????1??10?000111?) z |= 4'b1000; 
	if(x==?20'b11?????0?001??01111?) z |= 4'b1000; 
	if(x==?20'b111?1?11?110??0?1?1?) z |= 4'b1000; 
	if(x==?20'b?1??1?????00?1110?11) z |= 4'b1000; 
	if(x==?20'b?1?1??11?101010??1??) z |= 4'b0100; 
	if(x==?20'b?111???1010?01???11?) z |= 4'b0100; 
	if(x==?20'b1?1??1?0??0??1101?11) z |= 4'b1000; 
	if(x==?20'b?1?10?1??0??011?1?11) z |= 4'b0100; 
	if(x==?20'b?1??0?11111?0?0???01) z |= 4'b0100; 
	if(x==?20'b111???111110??0?1?1?) z |= 4'b1000; 
	if(x==?20'b1?1?11??101??010?1??) z |= 4'b1000; 
	if(x==?20'b?11111??0111?0??1?1?) z |= 4'b0100; 
	if(x==?20'b?1?????100?1110?1?11) z |= 4'b0100; 
	if(x==?20'b?1110??1?10?01???11?) z |= 4'b0100; 
	if(x==?20'b??1?11?0?111?0?0??01) z |= 4'b1000; 
	if(x==?20'b?1110??101??01???11?) z |= 4'b0100; 
	if(x==?20'b1???1?0?1110?00?1??1) z |= 4'b1000; 
	if(x==?20'b?1111????10?10??110?) z |= 4'b0100; 
	if(x==?20'b???10??1011?000?1??1) z |= 4'b0100; 
	if(x==?20'b111???10??0??101?1?1) z |= 4'b1000; 
	if(x==?20'b1???1??0?110?0001??1) z |= 4'b1000; 
	if(x==?20'b??1?0??1?0?1110?1?11) z |= 4'b0100; 
	if(x==?20'b??1?1???1?00?0111?11) z |= 4'b1000; 
	if(x==?20'b?1111???01??1?0?110?) z |= 4'b0100; 
	if(x==?20'b111?1????010??10?11?) z |= 4'b1000; 
	if(x==?20'b??1?1???1101?101?11?) z |= 4'b1000; 
	if(x==?20'b?1??1???1101?101?11?) z |= 4'b1000; 
	if(x==?20'b?11101???0??101??1?1) z |= 4'b0100; 
	if(x==?20'b???1?0?10111?00?1??1) z |= 4'b0100; 
	if(x==?20'b???111??000?00??1?11) z |= 4'b0100; 
	if(x==?20'b???101??000??1???101) z |= 4'b0100; 
	if(x==?20'b?11111??110??00?1?1?) z |= 4'b0100; 
	if(x==?20'b?1??1??01?0??0111?11) z |= 4'b1000; 
	if(x==?20'b111?1??0?01???10?11?) z |= 4'b1000; 
	if(x==?20'b???10?1?11??000?1?01) z |= 4'b0100; 
	if(x==?20'b???10?1?00??111???11) z |= 4'b0100; 
	if(x==?20'b1??????01110?0001??1) z |= 4'b1000; 
	if(x==?20'b?11?0?11???1111???11) z |= 4'b0100; 
	if(x==?20'b?11?11?01????111??11) z |= 4'b1000; 
	if(x==?20'b1?????11?000??001?11) z |= 4'b1000; 
	if(x==?20'b111?1??0??10??10?11?) z |= 4'b1000; 
	if(x==?20'b1?1???10100???0011??) z |= 4'b1000; 
	if(x==?20'b?11????1010?101??11?) z |= 4'b0100; 
	if(x==?20'b?????10?0111100?11??) z |= 4'b0100; 
	if(x==?20'b???10???0111000?1??1) z |= 4'b0100; 
	if(x==?20'b??1?1?001110??0?1??1) z |= 4'b1000; 
	if(x==?20'b??1????11011101??11?) z |= 4'b0100; 
	if(x==?20'b?1?????11011101??11?) z |= 4'b0100; 
	if(x==?20'b?????01?1110?00111??) z |= 4'b1000; 
	if(x==?20'b1?????10?000??1??101) z |= 4'b1000; 
	if(x==?20'b?11?1????010?101?11?) z |= 4'b1000; 
	if(x==?20'b?1??00?10111?0??1??1) z |= 4'b0100; 
	if(x==?20'b1????1?0??00?111??11) z |= 4'b1000; 
	if(x==?20'b111????1??10??01110?) z |= 4'b1000; 
	if(x==?20'b111???11?011?00?1?1?) z |= 4'b1000; 
	if(x==?20'b1????1?0??11?0001?01) z |= 4'b1000; 
	if(x==?20'b?1?10?11111???0???01) z |= 4'b0100; 
	if(x==?20'b?1?????0?001?100111?) z |= 4'b1000; 
	if(x==?20'b?1?10?1?011??11?1?1?) z |= 4'b0100; 
	if(x==?20'b1?1?11?0?111?0????01) z |= 4'b1000; 
	if(x==?20'b??1?0???100?001?111?) z |= 4'b0100; 
	if(x==?20'b??1?1?0?1110??001??1) z |= 4'b1000; 
	if(x==?20'b?111?1??101??10??10?) z |= 4'b0100; 
	if(x==?20'b1?1??1?0?110?11?1?1?) z |= 4'b1000; 
	if(x==?20'b?111?1??01?1?10??10?) z |= 4'b0100; 
	if(x==?20'b?1???0?1011100??1??1) z |= 4'b0100; 
	if(x==?20'b1?????101101??00?11?) z |= 4'b1000; 
	if(x==?20'b????001?100??1??110?) z |= 4'b0110; 
	if(x==?20'b?11????1?010?10?110?) z |= 4'b1000; 
	if(x==?20'b111???1??101?01??10?) z |= 4'b1000; 
	if(x==?20'b?1?1??11111?0?0???01) z |= 4'b0100; 
	if(x==?20'b??1101??010?00???11?) z |= 4'b0100; 
	if(x==?20'b111???1?1?10?01??10?) z |= 4'b1000; 
	if(x==?20'b???101??101100???11?) z |= 4'b0100; 
	if(x==?20'b?1111???0?11??1?110?) z |= 4'b0100; 
	if(x==?20'b1?1?11???111?0?0??01) z |= 4'b1000; 
	if(x==?20'b??1?1???1110?101?11?) z |= 4'b1000; 
	if(x==?20'b?1??1???1110?101?11?) z |= 4'b1000; 
	if(x==?20'b??11???1101?010??11?) z |= 4'b0100; 
	if(x==?20'b??1??1?01?0??1101?11) z |= 4'b1000; 
	if(x==?20'b?1???1??010?000??110) z |= 4'b0100; 
	if(x==?20'b?1?10?1??0??110?1?11) z |= 4'b0100; 
	if(x==?20'b11????10?010??00?11?) z |= 4'b1000; 
	if(x==?20'b?1?1???1010100??11??) z |= 4'b0100; 
	if(x==?20'b1?1?1???1010??0011??) z |= 4'b1000; 
	if(x==?20'b?11111??011??00?1?1?) z |= 4'b0100; 
	if(x==?20'b?1???1?01??0?1101?11) z |= 4'b1000; 
	if(x==?20'b??1????10111101??11?) z |= 4'b0100; 
	if(x==?20'b?1?????10111101??11?) z |= 4'b0100; 
	if(x==?20'b?1?10?1??11?011?1?1?) z |= 4'b0100; 
	if(x==?20'b11??1????101?010?11?) z |= 4'b1000; 
	if(x==?20'b1????1?01110?0?01??1) z |= 4'b1000; 
	if(x==?20'b1?1??1?0?11??1101?1?) z |= 4'b1000; 
	if(x==?20'b??1?0?1?0??1011?1?11) z |= 4'b0100; 
	if(x==?20'b?1??0?1??0?1011?1?11) z |= 4'b0100; 
	if(x==?20'b111???11?110?00?1?1?) z |= 4'b1000; 
	if(x==?20'b??1???1??010?000?110) z |= 4'b1000; 
	if(x==?20'b????110??001???1110?) z |= 4'b1000; 
	if(x==?20'b?????100?001??1?110?) z |= 4'b1001; 
	if(x==?20'b???10?1?01110?0?1??1) z |= 4'b0100; 
	if(x==?20'b?1??0?1?111?000???01) z |= 4'b0100; 
	if(x==?20'b????1??01110?0001??1) z |= 4'b1000; 
	if(x==?20'b??110???100??01?111?) z |= 4'b0100; 
	if(x==?20'b?1?10??1011?00??1??1) z |= 4'b0100; 
	if(x==?20'b1?1?1??0?110??001??1) z |= 4'b1000; 
	if(x==?20'b??1?1?1010?0?0?011??) z |= 4'b1000; 
	if(x==?20'b????0??10111000?1??1) z |= 4'b0100; 
	if(x==?20'b????1110?0?1?01011??) z |= 4'b1000; 
	if(x==?20'b1?1??1?0??0??0111?11) z |= 4'b1000; 
	if(x==?20'b??110??1111?000????1) z |= 4'b0100; 
	if(x==?20'b??1??1?0?111?000??01) z |= 4'b1000; 
	if(x==?20'b??1?1??01101?0?0?1?1) z |= 4'b1000; 
	if(x==?20'b?111???1?10?101??11?) z |= 4'b0100; 
	if(x==?20'b????01??0001?1???101) z |= 4'b0100; 
	if(x==?20'b?1?10?1?11??00??1?01) z |= 4'b0100; 
	if(x==?20'b11??1??0?111?000???1) z |= 4'b1000; 
	if(x==?20'b?111???101??101??11?) z |= 4'b0100; 
	if(x==?20'b?1??01?10?010?0?11??) z |= 4'b0100; 
	if(x==?20'b111?1????01??101?11?) z |= 4'b1000; 
	if(x==?20'b????0?1?00?1111???11) z |= 4'b0100; 
	if(x==?20'b11???????001?100111?) z |= 4'b1000; 
	if(x==?20'b1?????101110??00?11?) z |= 4'b1000; 
	if(x==?20'b??????101000??1??101) z |= 4'b1000; 
	if(x==?20'b111?1?????10?101?11?) z |= 4'b1000; 
	if(x==?20'b?1??00?1011??00?1??1) z |= 4'b0100; 
	if(x==?20'b??1?1?00?110?00?1??1) z |= 4'b1000; 
	if(x==?20'b??11????100?001?111?) z |= 4'b0100; 
	if(x==?20'b?????1?01?00?111??11) z |= 4'b1000; 
	if(x==?20'b?1??0??110110?0??1?1) z |= 4'b0100; 
	if(x==?20'b???101??011100???11?) z |= 4'b0100; 
	if(x==?20'b??11?10??001?00?11??) z |= 4'b0100; 
	if(x==?20'b??1?0??111??000?1?01) z |= 4'b0100; 
	if(x==?20'b??1?10011001????11??) z |= 4'b1100; 
	if(x==?20'b?1??10011001????11??) z |= 4'b1100; 
	if(x==?20'b?1111????10??10?110?) z |= 4'b0100; 
	if(x==?20'b1?1??1?0??11??001?01) z |= 4'b1000; 
	if(x==?20'b????0111?10?010?11??) z |= 4'b0100; 
	if(x==?20'b??1?0???100?100?111?) z |= 4'b0100; 
	if(x==?20'b?1??1??0??11?0001?01) z |= 4'b1000; 
	if(x==?20'b?1?10?1?111??00???01) z |= 4'b0100; 
	if(x==?20'b1???1??01110?00?1??1) z |= 4'b1000; 
	if(x==?20'b?1???0?1011?000?1??1) z |= 4'b0100; 
	if(x==?20'b??1?1?0??110?0001??1) z |= 4'b1000; 
	if(x==?20'b?1110??101?1?1???11?) z |= 4'b0100; 
	if(x==?20'b1?1??1??1?0??1101?11) z |= 4'b1000; 
	if(x==?20'b???10??10111?00?1??1) z |= 4'b0100; 
	if(x==?20'b1?1??1?0?111?00???01) z |= 4'b1000; 
	if(x==?20'b?1111???0?1??01?110?) z |= 4'b0100; 
	if(x==?20'b?1??00?1?11?000?1??1) z |= 4'b0100; 
	if(x==?20'b?11101???0??010??1?1) z |= 4'b0100; 
	if(x==?20'b???111??11??000?1?10) z |= 4'b0100; 
	if(x==?20'b111?1??01?10??1??11?) z |= 4'b1000; 
	if(x==?20'b111????1?01??01?110?) z |= 4'b1000; 
	if(x==?20'b?11??01?100???0011??) z |= 4'b1000; 
	if(x==?20'b?1?1??1??0?1011?1?11) z |= 4'b0100; 
	if(x==?20'b?1?????0?001?001111?) z |= 4'b1000; 
	if(x==?20'b111????1??10?01?110?) z |= 4'b1000; 
	if(x==?20'b1???1??0111??000??11) z |= 4'b1000; 
	if(x==?20'b?1???1??1110?1101?1?) z |= 4'b1000; 
	if(x==?20'b?1??00100100????11??) z |= 4'b1100; 
	if(x==?20'b111???10??0??010?1?1) z |= 4'b1000; 
	if(x==?20'b?111???1101?01???11?) z |= 4'b0100; 
	if(x==?20'b?1?1??1?111?000???01) z |= 4'b0100; 
	if(x==?20'b1?1??????100?100111?) z |= 4'b1000; 
	if(x==?20'b1???1???1110?0001??1) z |= 4'b1000; 
	if(x==?20'b?11????1010?010??11?) z |= 4'b0100; 
	if(x==?20'b??1???1?0111011?1?1?) z |= 4'b0100; 
	if(x==?20'b??1?0?1?1101?0??1?01) z |= 4'b0100; 
	if(x==?20'b??1????11011010??11?) z |= 4'b0100; 
	if(x==?20'b?1?????11011010??11?) z |= 4'b0100; 
	if(x==?20'b??1?1???1101?010?11?) z |= 4'b1000; 
	if(x==?20'b?1??1???1101?010?11?) z |= 4'b1000; 
	if(x==?20'b??1?1100110??0??1?1?) z |= 4'b1000; 
	if(x==?20'b?111???101?101???11?) z |= 4'b0100; 
	if(x==?20'b?1?10?11111?0?0????1) z |= 4'b0100; 
	if(x==?20'b??1?1100110???0?1?1?) z |= 4'b1000; 
	if(x==?20'b??11????001?010?111?) z |= 4'b0100; 
	if(x==?20'b?1?10?1??11?110?1?1?) z |= 4'b0100; 
	if(x==?20'b1?????11??11?0001?10) z |= 4'b1000; 
	if(x==?20'b??1?0?1?0??1110?1?11) z |= 4'b0100; 
	if(x==?20'b11?????0?10??100111?) z |= 4'b1000; 
	if(x==?20'b?1??0?1??0?1110?1?11) z |= 4'b0100; 
	if(x==?20'b???10??1?111000???11) z |= 4'b0100; 
	if(x==?20'b??1?01000010????11??) z |= 4'b1100; 
	if(x==?20'b???1???10111000?1??1) z |= 4'b0100; 
	if(x==?20'b1?1?11?0?111?0?0???1) z |= 4'b1000; 
	if(x==?20'b1?1??1???111?000??01) z |= 4'b1000; 
	if(x==?20'b111?1????101??10?11?) z |= 4'b1000; 
	if(x==?20'b1???1?11??00?0?01?11) z |= 4'b1000; 
	if(x==?20'b1?1??1?01110???01??1) z |= 4'b1000; 
	if(x==?20'b11???????100?010111?) z |= 4'b1000; 
	if(x==?20'b?1???1?01011??0?1?01) z |= 4'b1000; 
	if(x==?20'b111?1???1?10??10?11?) z |= 4'b1000; 
	if(x==?20'b???111?100??0?0?1?11) z |= 4'b0100; 
	if(x==?20'b???10?11?0??111???11) z |= 4'b0100; 
	if(x==?20'b?1?10?1?01110???1??1) z |= 4'b0100; 
	if(x==?20'b???1?1??0001?1???101) z |= 4'b0100; 
	if(x==?20'b?1?1????001?001?111?) z |= 4'b0100; 
	if(x==?20'b?1??1??01110?0?01??1) z |= 4'b1000; 
	if(x==?20'b?11?0?1?111?0?0???01) z |= 4'b0100; 
	if(x==?20'b??1?1??01110??001??1) z |= 4'b1000; 
	if(x==?20'b???1??1?00?1111???11) z |= 4'b0100; 
	if(x==?20'b?11?1????010?010?11?) z |= 4'b1000; 
	if(x==?20'b??1??1?01?0??0111?11) z |= 4'b1000; 
	if(x==?20'b1?????1?1000??1??101) z |= 4'b1000; 
	if(x==?20'b1?????111?00?0?01?11) z |= 4'b1000; 
	if(x==?20'b?1??0011?011?0??1?1?) z |= 4'b0100; 
	if(x==?20'b1???11?0??0??111??11) z |= 4'b1000; 
	if(x==?20'b?1??0011?011??0?1?1?) z |= 4'b0100; 
	if(x==?20'b??1???1?110100??1?01) z |= 4'b0100; 
	if(x==?20'b1????1??1?00?111??11) z |= 4'b1000; 
	if(x==?20'b111?1??0111??0?0???1) z |= 4'b1000; 
	if(x==?20'b????11??000?000?1?11) z |= 4'b0100; 
	if(x==?20'b?1??0??1011100??1??1) z |= 4'b0100; 
	if(x==?20'b??110????01?001?111?) z |= 4'b0100; 
	if(x==?20'b?1???1?01??0?0111?11) z |= 4'b1000; 
	if(x==?20'b??1?0??101110?0?1??1) z |= 4'b0100; 
	if(x==?20'b?11??1?0?111?0?0??01) z |= 4'b1000; 
	if(x==?20'b???111??00?10?0?1?11) z |= 4'b0100; 
	if(x==?20'b??????11?000?0001?11) z |= 4'b1000; 
	if(x==?20'b?11?1????101?101?11?) z |= 4'b1000; 
	if(x==?20'b1?1??1?0?11??0111?1?) z |= 4'b1000; 
	if(x==?20'b?111011??1??101??1??) z |= 4'b0100; 
	if(x==?20'b?11????1101?101??11?) z |= 4'b0100; 
	if(x==?20'b?1???1??1011??001?01) z |= 4'b1000; 
	if(x==?20'b?????011100???1?110?) z |= 4'b0100; 
	if(x==?20'b1??????011?0?0001?11) z |= 4'b1000; 
	if(x==?20'b?11??11011???1101???) z |= 4'b1000; 
	if(x==?20'b111??110??1??101?1??) z |= 4'b1000; 
	if(x==?20'b?1110??1?1110?0????1) z |= 4'b0100; 
	if(x==?20'b??1????01101?000?1?1) z |= 4'b1000; 
	if(x==?20'b?111???1010??10??11?) z |= 4'b0100; 
	if(x==?20'b???10???0?11000?1?11) z |= 4'b0100; 
	if(x==?20'b111????1??01?10011??) z |= 4'b1000; 
	if(x==?20'b?1111???10??001?11??) z |= 4'b0100; 
	if(x==?20'b?1??0???1011000??1?1) z |= 4'b0100; 
	if(x==?20'b?11?011???11011?1???) z |= 4'b0100; 
	if(x==?20'b??1????10111010??11?) z |= 4'b0100; 
	if(x==?20'b?1?????10111010??11?) z |= 4'b0100; 
	if(x==?20'b????11?0?001???1110?) z |= 4'b1000; 
	if(x==?20'b?1110??1?10??10??11?) z |= 4'b0100; 
	if(x==?20'b??1?1???1110?010?11?) z |= 4'b1000; 
	if(x==?20'b?1??1???1110?010?11?) z |= 4'b1000; 
	if(x==?20'b?1110??101???10??11?) z |= 4'b0100; 
	if(x==?20'b?11100?111???0??1??1) z |= 4'b0100; 
	if(x==?20'b1?1?1??01110??0?1??1) z |= 4'b1000; 
	if(x==?20'b111?1????010?01??11?) z |= 4'b1000; 
	if(x==?20'b??????101101?000?11?) z |= 4'b1000; 
	if(x==?20'b???111??000??00?1?11) z |= 4'b0100; 
	if(x==?20'b?11?1???01?1?01?110?) z |= 4'b0100; 
	if(x==?20'b?1?10??10111?0??1??1) z |= 4'b0100; 
	if(x==?20'b11?????0??01?001111?) z |= 4'b1000; 
	if(x==?20'b??1101??101?00???11?) z |= 4'b0100; 
	if(x==?20'b111?1??0?01??01??11?) z |= 4'b1000; 
	if(x==?20'b11????10?101??00?11?) z |= 4'b1000; 
	if(x==?20'b?1?1??1??0?1110?1?11) z |= 4'b0100; 
	if(x==?20'b1?????11?000?00?1?11) z |= 4'b1000; 
	if(x==?20'b????01??1011000??11?) z |= 4'b0100; 
	if(x==?20'b111?1?00??11??0?1??1) z |= 4'b1000; 
	if(x==?20'b111?1??0??10?01??11?) z |= 4'b1000; 
	if(x==?20'b?111???1?10?010??11?) z |= 4'b0100; 
	if(x==?20'b?11????0?001??01111?) z |= 4'b1000; 
	if(x==?20'b11??1??0111??0?0??11) z |= 4'b1000; 
	if(x==?20'b?111???101??010??11?) z |= 4'b0100; 
	if(x==?20'b??1???1?0111110?1?1?) z |= 4'b0100; 
	if(x==?20'b1?1?1??0111???00??11) z |= 4'b1000; 
	if(x==?20'b111????01?0??000??11) z |= 4'b1000; 
	if(x==?20'b?111?0?111??00??1??1) z |= 4'b0100; 
	if(x==?20'b1?1?1???1110??001??1) z |= 4'b1000; 
	if(x==?20'b1?1??1??1?0??0111?11) z |= 4'b1000; 
	if(x==?20'b?1?101???001?00?11??) z |= 4'b0100; 
	if(x==?20'b????1?111?00?0?01?11) z |= 4'b1000; 
	if(x==?20'b111????01??0?000??11) z |= 4'b1000; 
	if(x==?20'b??1?????0011010?111?) z |= 4'b0100; 
	if(x==?20'b?1?10?1?011?0?0?1??1) z |= 4'b0100; 
	if(x==?20'b?1?10??1?11100????11) z |= 4'b0100; 
	if(x==?20'b?1?1???1011100??1??1) z |= 4'b0100; 
	if(x==?20'b????1?11101?01??01??) z |= 4'b0100; 
	if(x==?20'b??110??1?1110?0???11) z |= 4'b0100; 
	if(x==?20'b111?1????01??010?11?) z |= 4'b1000; 
	if(x==?20'b?1110???0??1000???11) z |= 4'b0100; 
	if(x==?20'b?1110????0?1000???11) z |= 4'b0100; 
	if(x==?20'b?1?10?1?111?000????1) z |= 4'b0100; 
	if(x==?20'b1?1??1?0?110?0?01??1) z |= 4'b1000; 
	if(x==?20'b?1?1????001?100?111?) z |= 4'b0100; 
	if(x==?20'b111??????100??10111?) z |= 4'b1000; 
	if(x==?20'b111?1?0???11??001??1) z |= 4'b1000; 
	if(x==?20'b111?1?????10?010?11?) z |= 4'b1000; 
	if(x==?20'b????11?01?0??111??11) z |= 4'b1000; 
	if(x==?20'b??1?1?0?1110?00?1??1) z |= 4'b1000; 
	if(x==?20'b????11?100?10?0?1?11) z |= 4'b0100; 
	if(x==?20'b?1???1??1110?0111?1?) z |= 4'b1000; 
	if(x==?20'b????0?11?0?1111???11) z |= 4'b0100; 
	if(x==?20'b?111????001?0?1?111?) z |= 4'b0100; 
	if(x==?20'b111??11?11???1101???) z |= 4'b1000; 
	if(x==?20'b?1??0??1011?000?1??1) z |= 4'b0100; 
	if(x==?20'b??1?1??0?110?0001??1) z |= 4'b1000; 
	if(x==?20'b1?1??????100?001111?) z |= 4'b1000; 
	if(x==?20'b1?1??1?0?111?000???1) z |= 4'b1000; 
	if(x==?20'b1?????11??00?0001?11) z |= 4'b1000; 
	if(x==?20'b1?????101101?00??11?) z |= 4'b1000; 
	if(x==?20'b??110????01?100?111?) z |= 4'b0100; 
	if(x==?20'b11??????1?01?100111?) z |= 4'b1000; 
	if(x==?20'b????11?1?101??1001??) z |= 4'b1000; 
	if(x==?20'b?1???0?10111?00?1??1) z |= 4'b0100; 
	if(x==?20'b?1??11??000?00??1?11) z |= 4'b0100; 
	if(x==?20'b1?????111110??001?1?) z |= 4'b1000; 
	if(x==?20'b?1??01??000??1???101) z |= 4'b0100; 
	if(x==?20'b????11?11?10??1001??) z |= 4'b1000; 
	if(x==?20'b???111??011100??1?1?) z |= 4'b0100; 
	if(x==?20'b?1??0?1?11??000?1?01) z |= 4'b0100; 
	if(x==?20'b??1????01110?0001??1) z |= 4'b1000; 
	if(x==?20'b?1??0?1?00??111???11) z |= 4'b0100; 
	if(x==?20'b?1?????01110?0001??1) z |= 4'b1000; 
	if(x==?20'b??1?111?111?00????10) z |= 4'b0100; 
	if(x==?20'b???10?1?11?1000?1??1) z |= 4'b0100; 
	if(x==?20'b??1101??010??00??11?) z |= 4'b0100; 
	if(x==?20'b??1???11?000??001?11) z |= 4'b1000; 
	if(x==?20'b??????101110?000?11?) z |= 4'b1000; 
	if(x==?20'b?111?11???11011?1???) z |= 4'b0100; 
	if(x==?20'b???101??1011?00??11?) z |= 4'b0100; 
	if(x==?20'b??1?0???0111000?1??1) z |= 4'b0100; 
	if(x==?20'b?1??0???0111000?1??1) z |= 4'b0100; 
	if(x==?20'b1?1?????1100?10?111?) z |= 4'b1000; 
	if(x==?20'b111????0111??000???1) z |= 4'b1000; 
	if(x==?20'b1????1?01?11?0001??1) z |= 4'b1000; 
	if(x==?20'b????01??0111000??11?) z |= 4'b0100; 
	if(x==?20'b??1???10?000??1??101) z |= 4'b1000; 
	if(x==?20'b11????10?010?00??11?) z |= 4'b1000; 
	if(x==?20'b1?1?1???1010?00?11??) z |= 4'b1000; 
	if(x==?20'b111?111???11??111???) z |= 4'b1000; 
	if(x==?20'b??1??1?0??00?111??11) z |= 4'b1000; 
	if(x==?20'b?1?1???10101?00?11??) z |= 4'b0100; 
	if(x==?20'b?1???111?111??00??10) z |= 4'b1000; 
	if(x==?20'b?1110????111000????1) z |= 4'b0100; 
	if(x==?20'b??1??1?0??11?0001?01) z |= 4'b1000; 
	if(x==?20'b?1111???10??100?11??) z |= 4'b0100; 
	if(x==?20'b?11?01100??0?00?1?1?) z |= 4'b1100; 
	if(x==?20'b?1?1????0011?01?111?) z |= 4'b0100; 
	if(x==?20'b?1?10??1011??00?1??1) z |= 4'b0100; 
	if(x==?20'b1?1?1??0?110?00?1??1) z |= 4'b1000; 
	if(x==?20'b??1???101101??00?11?) z |= 4'b1000; 
	if(x==?20'b?1????101101??00?11?) z |= 4'b1000; 
	if(x==?20'b1???1?0?100???0011??) z |= 4'b1000; 
	if(x==?20'b111????1??01?00111??) z |= 4'b1000; 
	if(x==?20'b?11?01??010?00???11?) z |= 4'b0100; 
	if(x==?20'b?1?10?1?11???00?1?01) z |= 4'b0100; 
	if(x==?20'b??1?01??101100???11?) z |= 4'b0100; 
	if(x==?20'b??11111?111??0????10) z |= 4'b0100; 
	if(x==?20'b?1??01??101100???11?) z |= 4'b0100; 
	if(x==?20'b????0?11100???1?110?) z |= 4'b0100; 
	if(x==?20'b1?????101110?00??11?) z |= 4'b1000; 
	if(x==?20'b???1?0?1?00100??11??) z |= 4'b0100; 
	if(x==?20'b?111011??1??010??1??) z |= 4'b0100; 
	if(x==?20'b?11????1101?010??11?) z |= 4'b0100; 
	if(x==?20'b1???1?111?0???001?11) z |= 4'b1000; 
	if(x==?20'b1???11??1?0??111??11) z |= 4'b1000; 
	if(x==?20'b???1??11?0?1111???11) z |= 4'b0100; 
	if(x==?20'b??1?111?00??111????1) z |= 4'b0100; 
	if(x==?20'b?11???10?010??00?11?) z |= 4'b1000; 
	if(x==?20'b???101??0111?00??11?) z |= 4'b0100; 
	if(x==?20'b?1?1???1011?000?1??1) z |= 4'b0100; 
	if(x==?20'b1?1?1????110?0001??1) z |= 4'b1000; 
	if(x==?20'b11???111?111??0???10) z |= 4'b1000; 
	if(x==?20'b?11?1????101?010?11?) z |= 4'b1000; 
	if(x==?20'b??1??1?01110?0?01??1) z |= 4'b1000; 
	if(x==?20'b1?1??1?0??11?00?1?01) z |= 4'b1000; 
	if(x==?20'b11?????0111??000??11) z |= 4'b1000; 
	if(x==?20'b???111?1?0?100??1?11) z |= 4'b0100; 
	if(x==?20'b?1??0?1?01110?0?1??1) z |= 4'b0100; 
	if(x==?20'b?1?1??1?11??000?1?01) z |= 4'b0100; 
	if(x==?20'b111??110??1??010?1??) z |= 4'b1000; 
	if(x==?20'b??11?????011001?111?) z |= 4'b0100; 
	if(x==?20'b?1?1??1?00??111???11) z |= 4'b0100; 
	if(x==?20'b????0011010???1?11??) z |= 4'b0100; 
	if(x==?20'b??????11100?0?1?110?) z |= 4'b0100; 
	if(x==?20'b?11?0???100??01?111?) z |= 4'b0100; 
	if(x==?20'b?1???111??00?111???1) z |= 4'b1000; 
	if(x==?20'b??110????111000???11) z |= 4'b0100; 
	if(x==?20'b???110?11001????11??) z |= 4'b0100; 
	if(x==?20'b1???1?011001????11??) z |= 4'b1000; 
	if(x==?20'b????11???001??10110?) z |= 4'b1000; 
	if(x==?20'b??110?1??0??111???11) z |= 4'b0100; 
	if(x==?20'b1?1????1?100???1110?) z |= 4'b1000; 
	if(x==?20'b?11?0??1111?000????1) z |= 4'b0100; 
	if(x==?20'b????1100?010??1?11??) z |= 4'b1000; 
	if(x==?20'b1?1???11??00??001?11) z |= 4'b1000; 
	if(x==?20'b1?1??1????00?111??11) z |= 4'b1000; 
	if(x==?20'b1?1??1????11?0001?01) z |= 4'b1000; 
	if(x==?20'b?11?1??0?111?000???1) z |= 4'b1000; 
	if(x==?20'b?1?10?1?11?100??1??1) z |= 4'b0100; 
	if(x==?20'b11???1?0??0??111??11) z |= 4'b1000; 
	if(x==?20'b??1???101110??00?11?) z |= 4'b1000; 
	if(x==?20'b?1????101110??00?11?) z |= 4'b1000; 
	if(x==?20'b?111???1101??10??11?) z |= 4'b0100; 
	if(x==?20'b1?1??1?01?11??001??1) z |= 4'b1000; 
	if(x==?20'b???1011111??0?0?1?1?) z |= 4'b0100; 
	if(x==?20'b??1?01??011100???11?) z |= 4'b0100; 
	if(x==?20'b?1??01??011100???11?) z |= 4'b0100; 
	if(x==?20'b?1110??111??00??1??1) z |= 4'b0100; 
	if(x==?20'b???10??100??01???111) z |= 4'b0100; 
	if(x==?20'b?111???101?1?10??11?) z |= 4'b0100; 
	if(x==?20'b?11??10??001?00?11??) z |= 4'b0100; 
	if(x==?20'b??1?0??111?1000?1??1) z |= 4'b0100; 
	if(x==?20'b?????11?101?101?01??) z |= 4'b0100; 
	if(x==?20'b?????11??101?10101??) z |= 4'b1000; 
	if(x==?20'b?1??1??01?11?0001??1) z |= 4'b1000; 
	if(x==?20'b11??????1?01?001111?) z |= 4'b1000; 
	if(x==?20'b11????1?1101??00?11?) z |= 4'b1000; 
	if(x==?20'b111?1????101?01??11?) z |= 4'b1000; 
	if(x==?20'b1?1??1?01110?0??1??1) z |= 4'b1000; 
	if(x==?20'b?1?????11100?0?0111?) z |= 4'b1000; 
	if(x==?20'b?111?11111???11?1???) z |= 4'b0100; 
	if(x==?20'b1???1110??11?0?01?1?) z |= 4'b1000; 
	if(x==?20'b111?1???1?10?01??11?) z |= 4'b1000; 
	if(x==?20'b1???1??0??00??10?111) z |= 4'b1000; 
	if(x==?20'b111?1??0??11??001??1) z |= 4'b1000; 
	if(x==?20'b?111?1??010?00???11?) z |= 4'b0100; 
	if(x==?20'b?1?10?1?0111??0?1??1) z |= 4'b0100; 
	if(x==?20'b??11?1??101100???11?) z |= 4'b0100; 
	if(x==?20'b??1?1??01110?00?1??1) z |= 4'b1000; 
	if(x==?20'b????0111101??1??01??) z |= 4'b0100; 
	if(x==?20'b????011101?1?1??01??) z |= 4'b0100; 
	if(x==?20'b?????10011?0??1011??) z |= 4'b1000; 
	if(x==?20'b??1???1?1101?00?1?01) z |= 4'b0100; 
	if(x==?20'b?11101???10?00???11?) z |= 4'b0100; 
	if(x==?20'b111???1??010??00?11?) z |= 4'b1000; 
	if(x==?20'b?1??0??10111?00?1??1) z |= 4'b0100; 
	if(x==?20'b11??1?0?100????011??) z |= 4'b1000; 
	if(x==?20'b1?1??1?0111??0?0??11) z |= 4'b1000; 
	if(x==?20'b?11101??01??00???11?) z |= 4'b0100; 
	if(x==?20'b????1110?101??1?01??) z |= 4'b1000; 
	if(x==?20'b??1?11??11??000?1?10) z |= 4'b0100; 
	if(x==?20'b?1??11??11??000?1?10) z |= 4'b0100; 
	if(x==?20'b????001?0?110?1?11??) z |= 4'b0100; 
	if(x==?20'b1?1??1??1110?0?01??1) z |= 4'b1000; 
	if(x==?20'b????11101?10??1?01??) z |= 4'b1000; 
	if(x==?20'b?1???1??1011?00?1?01) z |= 4'b1000; 
	if(x==?20'b111???10?01???00?11?) z |= 4'b1000; 
	if(x==?20'b????1??0??00?101?111) z |= 4'b1000; 
	if(x==?20'b??1?1??0111??000??11) z |= 4'b1000; 
	if(x==?20'b?1?10?1??1110?0???11) z |= 4'b0100; 
	if(x==?20'b?1?1??1?01110?0?1??1) z |= 4'b0100; 
	if(x==?20'b????0??100??101??111) z |= 4'b0100; 
	if(x==?20'b111???10??10??00?11?) z |= 4'b1000; 
	if(x==?20'b??1?1???100?000?111?) z |= 4'b0100; 
	if(x==?20'b??11?0?1?0010???11??) z |= 4'b0100; 
	if(x==?20'b??1?1???1110?0001??1) z |= 4'b1000; 
	if(x==?20'b???10??101?101???11?) z |= 4'b0100; 
	if(x==?20'b1???1?11??0??0001?11) z |= 4'b1000; 
	if(x==?20'b?11?????001?010?111?) z |= 4'b0100; 
	if(x==?20'b?????11101?101??01??) z |= 4'b0100; 
	if(x==?20'b???111?1?0??000?1?11) z |= 4'b0100; 
	if(x==?20'b??1???11??11?0001?10) z |= 4'b1000; 
	if(x==?20'b?1????11??11?0001?10) z |= 4'b1000; 
	if(x==?20'b?11????0?10??100111?) z |= 4'b1000; 
	if(x==?20'b?1??0??1?111000???11) z |= 4'b0100; 
	if(x==?20'b?1?????10111000?1??1) z |= 4'b0100; 
	if(x==?20'b1?1??1111??0?0?0??11) z |= 4'b1000; 
	if(x==?20'b1???1??01?10??10?11?) z |= 4'b1000; 
	if(x==?20'b1?????111?0??0001?11) z |= 4'b1000; 
	if(x==?20'b??1?1?11??00?0?01?11) z |= 4'b1000; 
	if(x==?20'b?1?????1?001?000111?) z |= 4'b1000; 
	if(x==?20'b?11??????100?010111?) z |= 4'b1000; 
	if(x==?20'b??11?????011100?111?) z |= 4'b0100; 
	if(x==?20'b?1??11?100??0?0?1?11) z |= 4'b0100; 
	if(x==?20'b?1?1111?0??10?0???11) z |= 4'b0100; 
	if(x==?20'b??1?0?110???111???11) z |= 4'b0100; 
	if(x==?20'b?1??0?11?0??111???11) z |= 4'b0100; 
	if(x==?20'b?1???1??0001?1???101) z |= 4'b0100; 
	if(x==?20'b?1????1?00?1111???11) z |= 4'b0100; 
	if(x==?20'b??1???1?1000??1??101) z |= 4'b1000; 
	if(x==?20'b??1???111?00?0?01?11) z |= 4'b1000; 
	if(x==?20'b?1????111?00?0?01?11) z |= 4'b1000; 
	if(x==?20'b??1?11?0??0??111??11) z |= 4'b1000; 
	if(x==?20'b???111???0?1000?1?11) z |= 4'b0100; 
	if(x==?20'b????0?1?100??01?110?) z |= 4'b0110; 
	if(x==?20'b??1??1??1?00?111??11) z |= 4'b1000; 
	if(x==?20'b??????111110?0001?1?) z |= 4'b1000; 
	if(x==?20'b??????1?100?001?110?) z |= 4'b0100; 
	if(x==?20'b?11?0????01?001?111?) z |= 4'b0100; 
	if(x==?20'b?1?10?1?11??000?1??1) z |= 4'b0100; 
	if(x==?20'b?1??11?0???0?111??11) z |= 4'b1000; 
	if(x==?20'b????11??0111000?1?1?) z |= 4'b0100; 
	if(x==?20'b??1?11??00?10?0?1?11) z |= 4'b0100; 
	if(x==?20'b?1??11??00?10?0?1?11) z |= 4'b0100; 
	if(x==?20'b11????10?101?00??11?) z |= 4'b1000; 
	if(x==?20'b??1?0?1??0?1111???11) z |= 4'b0100; 
	if(x==?20'b??1101??101??00??11?) z |= 4'b0100; 
	if(x==?20'b111?1?1?1??0?0?0??11) z |= 4'b1000; 
	if(x==?20'b?1???1?01?0??111??11) z |= 4'b1000; 
	if(x==?20'b????11???001?0?1110?) z |= 4'b1000; 
	if(x==?20'b??1????011?0?0001?11) z |= 4'b1000; 
	if(x==?20'b?1110?1?11?10???1??1) z |= 4'b0100; 
	if(x==?20'b?11?????100?100?111?) z |= 4'b0100; 
	if(x==?20'b1?1?1??0111??00???11) z |= 4'b1000; 
	if(x==?20'b??111???100??00?111?) z |= 4'b0100; 
	if(x==?20'b1?1?1???1110?00?1??1) z |= 4'b1000; 
	if(x==?20'b?????1???001?100110?) z |= 4'b1001; 
	if(x==?20'b111??1?01?11???01??1) z |= 4'b1000; 
	if(x==?20'b?111?1?10??10?0???11) z |= 4'b0100; 
	if(x==?20'b?111?0?111???00?1??1) z |= 4'b0100; 
	if(x==?20'b1?1??1?0??11?0001??1) z |= 4'b1000; 
	if(x==?20'b?1??0???0?11000?1?11) z |= 4'b0100; 
	if(x==?20'b?1?11???001??1??110?) z |= 4'b0100; 
	if(x==?20'b?111????001??10?111?) z |= 4'b0100; 
	if(x==?20'b?1?10??1?111?00???11) z |= 4'b0100; 
	if(x==?20'b?1?1???10111?00?1??1) z |= 4'b0100; 
	if(x==?20'b????1?11101??10?01??) z |= 4'b0100; 
	if(x==?20'b?1110???11??000?1??1) z |= 4'b0100; 
	if(x==?20'b11?????1?001?00?111?) z |= 4'b1000; 
	if(x==?20'b111??????100?01?111?) z |= 4'b1000; 
	if(x==?20'b111?1?0???11?00?1??1) z |= 4'b1000; 
	if(x==?20'b1?1????1?100??1?110?) z |= 4'b1000; 
	if(x==?20'b?11??????001?001111?) z |= 4'b1000; 
	if(x==?20'b1???1?????00?101?111) z |= 4'b1000; 
	if(x==?20'b?1?11???001???1?110?) z |= 4'b0100; 
	if(x==?20'b1?1?1???111??000??11) z |= 4'b1000; 
	if(x==?20'b???1???100??101??111) z |= 4'b0100; 
	if(x==?20'b????11?1?101?01?01??) z |= 4'b1000; 
	if(x==?20'b???111??0?1?000?1?11) z |= 4'b0100; 
	if(x==?20'b1?????111110?00?1?1?) z |= 4'b1000; 
	if(x==?20'b111????0??11?0001??1) z |= 4'b1000; 
	if(x==?20'b?1??11??000??00?1?11) z |= 4'b0100; 
	if(x==?20'b????11?11?10?01?01??) z |= 4'b1000; 
	if(x==?20'b?11????0??01?001111?) z |= 4'b1000; 
	if(x==?20'b?1110?????0?000?1?11) z |= 4'b0100; 
	if(x==?20'b?11?01??101?00???11?) z |= 4'b0100; 
	if(x==?20'b?11???10?101??00?11?) z |= 4'b1000; 
	if(x==?20'b???111??0111?00?1?1?) z |= 4'b0100; 
	if(x==?20'b????0?1?00??011?1?11) z |= 4'b0100; 
	if(x==?20'b?1?1???1?111000???11) z |= 4'b0100; 
	if(x==?20'b??1???11?000?00?1?11) z |= 4'b1000; 
	if(x==?20'b?????1?0??00?1101?11) z |= 4'b1000; 
	if(x==?20'b????1?111?0??0001?11) z |= 4'b1000; 
	if(x==?20'b??111???10??000?111?) z |= 4'b0100; 
	if(x==?20'b?11?1??0111??0?0??11) z |= 4'b1000; 
	if(x==?20'b??11??110???111???11) z |= 4'b0100; 
	if(x==?20'b????0?11010?0?1?11??) z |= 4'b0100; 
	if(x==?20'b?1?1??11?0??111???11) z |= 4'b0100; 
	if(x==?20'b??11??1?010101???1??) z |= 4'b0100; 
	if(x==?20'b?11?1???100?00??111?) z |= 4'b0100; 
	if(x==?20'b???1???1001?010?11??) z |= 4'b0100; 
	if(x==?20'b1??????01??0?101?111) z |= 4'b1000; 
	if(x==?20'b1?1?1?11??0???001?11) z |= 4'b1000; 
	if(x==?20'b1?1?11????0??111??11) z |= 4'b1000; 
	if(x==?20'b1?1?111?111??0?0??1?) z |= 4'b1000; 
	if(x==?20'b1???1????100?01011??) z |= 4'b1000; 
	if(x==?20'b11?????1??01?000111?) z |= 4'b1000; 
	if(x==?20'b?1?111?1?0??00??1?11) z |= 4'b0100; 
	if(x==?20'b???10???0??1101??111) z |= 4'b0100; 
	if(x==?20'b????011101??101??1??) z |= 4'b0100; 
	if(x==?20'b????11?0?010??1011??) z |= 4'b1000; 
	if(x==?20'b?1110??111?1?0??1??1) z |= 4'b0100; 
	if(x==?20'b????11?1?0?1000?1?11) z |= 4'b0100; 
	if(x==?20'b?11?0??1?1110?0???11) z |= 4'b0100; 
	if(x==?20'b11??11?????0?111??11) z |= 4'b1000; 
	if(x==?20'b?????11?101?010?01??) z |= 4'b0100; 
	if(x==?20'b111?1??01?11??0?1??1) z |= 4'b1000; 
	if(x==?20'b??11??1??0?1111???11) z |= 4'b0100; 
	if(x==?20'b11???1??1?0??111??11) z |= 4'b1000; 
	if(x==?20'b11???1??1010??10?1??) z |= 4'b1000; 
	if(x==?20'b1?1?????11?0?0001?11) z |= 4'b1000; 
	if(x==?20'b?1?1?111?1110?0???1?) z |= 4'b0100; 
	if(x==?20'b?????11??101?01001??) z |= 4'b1000; 
	if(x==?20'b??1???11??00?0001?11) z |= 4'b1000; 
	if(x==?20'b??1???101101?00??11?) z |= 4'b1000; 
	if(x==?20'b?1????101101?00??11?) z |= 4'b1000; 
	if(x==?20'b?11?0????01?100?111?) z |= 4'b0100; 
	if(x==?20'b???10??11?1?101??11?) z |= 4'b0100; 
	if(x==?20'b1?1????011???0001?11) z |= 4'b1000; 
	if(x==?20'b1???1??0?1?1?101?11?) z |= 4'b1000; 
	if(x==?20'b??1???111110??001?1?) z |= 4'b1000; 
	if(x==?20'b?1????111110??001?1?) z |= 4'b1000; 
	if(x==?20'b?1??1??0??00??111?11) z |= 4'b1000; 
	if(x==?20'b1???1?0?1?00?00?11??) z |= 4'b1000; 
	if(x==?20'b?1?1????0?11000?1?11) z |= 4'b0100; 
	if(x==?20'b??1?11??011100??1?1?) z |= 4'b0100; 
	if(x==?20'b?1??11??011100??1?1?) z |= 4'b0100; 
	if(x==?20'b?1110?1?11??0?0?1??1) z |= 4'b0100; 
	if(x==?20'b?111???111?100??1??1) z |= 4'b0100; 
	if(x==?20'b?1??0?1?11?1000?1??1) z |= 4'b0100; 
	if(x==?20'b?11?01??010??00??11?) z |= 4'b0100; 
	if(x==?20'b111?1???1?11??001??1) z |= 4'b1000; 
	if(x==?20'b??1?01??1011?00??11?) z |= 4'b0100; 
	if(x==?20'b?1??01??1011?00??11?) z |= 4'b0100; 
	if(x==?20'b???1?0?1?001?00?11??) z |= 4'b0100; 
	if(x==?20'b1???1?111?0??00?1?11) z |= 4'b1000; 
	if(x==?20'b??1??1?01?11?0001??1) z |= 4'b1000; 
	if(x==?20'b?1?10?????11000?1?11) z |= 4'b0100; 
	if(x==?20'b??????1?100?100?110?) z |= 4'b0110; 
	if(x==?20'b????0??100??010??111) z |= 4'b0100; 
	if(x==?20'b?11???10?010?00??11?) z |= 4'b1000; 
	if(x==?20'b111???1?1??0?000??11) z |= 4'b1000; 
	if(x==?20'b111??1?0??11?0?01??1) z |= 4'b1000; 
	if(x==?20'b??????11100??10?110?) z |= 4'b0100; 
	if(x==?20'b?????1???001?001110?) z |= 4'b1000; 
	if(x==?20'b?11?1???00??000?1?11) z |= 4'b0100; 
	if(x==?20'b??1?011111?10???1?1?) z |= 4'b0100; 
	if(x==?20'b?1??11101?11???01?1?) z |= 4'b1000; 
	if(x==?20'b?111?1??0??1000???11) z |= 4'b0100; 
	if(x==?20'b????1??0??00?010?111) z |= 4'b1000; 
	if(x==?20'b???111?1?0?1?00?1?11) z |= 4'b0100; 
	if(x==?20'b?111?1??101?00???11?) z |= 4'b0100; 
	if(x==?20'b111???1??101??00?11?) z |= 4'b1000; 
	if(x==?20'b???1??1?00??011?1?11) z |= 4'b0100; 
	if(x==?20'b111????1?001??0?111?) z |= 4'b1000; 
	if(x==?20'b111???1?1?10??00?11?) z |= 4'b1000; 
	if(x==?20'b?111?1??01?100???11?) z |= 4'b0100; 
	if(x==?20'b1????1????00?1101?11) z |= 4'b1000; 
	if(x==?20'b?1??1?0?100??0?011??) z |= 4'b1000; 
	if(x==?20'b??1?1?0?100???0011??) z |= 4'b1000; 
	if(x==?20'b1?1???11??00?00?1?11) z |= 4'b1000; 
	if(x==?20'b????0?11111?00????01) z |= 4'b0100; 
	if(x==?20'b?1?111??0?1?00??1?11) z |= 4'b0100; 
	if(x==?20'b????0?1?00??110?1?11) z |= 4'b0100; 
	if(x==?20'b11??1100???0???01?1?) z |= 4'b1000; 
	if(x==?20'b?11?111?111??0????10) z |= 4'b0100; 
	if(x==?20'b?1?10?1?11?1?00?1??1) z |= 4'b0100; 
	if(x==?20'b????11?0?111??00??01) z |= 4'b1000; 
	if(x==?20'b??1???101110?00??11?) z |= 4'b1000; 
	if(x==?20'b?1????101110?00??11?) z |= 4'b1000; 
	if(x==?20'b?1???0?1?00100??11??) z |= 4'b0100; 
	if(x==?20'b?1??1?111?0??0?01?11) z |= 4'b1000; 
	if(x==?20'b??1??0?1?0010?0?11??) z |= 4'b0100; 
	if(x==?20'b??1?1?111?0???001?11) z |= 4'b1000; 
	if(x==?20'b??1?11??1?0??111??11) z |= 4'b1000; 
	if(x==?20'b1?1??1?01?11?00?1??1) z |= 4'b1000; 
	if(x==?20'b??1???110??1111???11) z |= 4'b0100; 
	if(x==?20'b?1????11?0?1111???11) z |= 4'b0100; 
	if(x==?20'b??1?01??0111?00??11?) z |= 4'b0100; 
	if(x==?20'b?1??01??0111?00??11?) z |= 4'b0100; 
	if(x==?20'b?1110??111???00?1??1) z |= 4'b0100; 
	if(x==?20'b?1?1?01?0101?0???1??) z |= 4'b0100; 
	if(x==?20'b????0?1101??101??11?) z |= 4'b0100; 
	if(x==?20'b???10??100???10??111) z |= 4'b0100; 
	if(x==?20'b?1??1?111??0??001?11) z |= 4'b1000; 
	if(x==?20'b?1??11??1??0?111??11) z |= 4'b1000; 
	if(x==?20'b?11??111?111??0???10) z |= 4'b1000; 
	if(x==?20'b??111????01?10??110?) z |= 4'b0100; 
	if(x==?20'b1?1?1?11?11???001?1?) z |= 4'b1000; 
	if(x==?20'b11????1?1101?00??11?) z |= 4'b1000; 
	if(x==?20'b?1?111?1?11?00??1?1?) z |= 4'b0100; 
	if(x==?20'b1?1??10?1010??0??1??) z |= 4'b1000; 
	if(x==?20'b?11????0111??000??11) z |= 4'b1000; 
	if(x==?20'b??1?11?10??100??1?11) z |= 4'b0100; 
	if(x==?20'b?????10011?0?10?11??) z |= 4'b1000; 
	if(x==?20'b?1??11?1?0?100??1?11) z |= 4'b0100; 
	if(x==?20'b????11?0??10?101?11?) z |= 4'b1000; 
	if(x==?20'b??1?11?1?0?10?0?1?11) z |= 4'b0100; 
	if(x==?20'b??111?1?01??101??1??) z |= 4'b0100; 
	if(x==?20'b1???1??0??00?01??111) z |= 4'b1000; 
	if(x==?20'b111?1??0??11?00?1??1) z |= 4'b1000; 
	if(x==?20'b?11??????011001?111?) z |= 4'b0100; 
	if(x==?20'b?1?1??1?11?1000?1??1) z |= 4'b0100; 
	if(x==?20'b?????1?0??00?0111?11) z |= 4'b1000; 
	if(x==?20'b1???1??0?101??00?1?1) z |= 4'b1000; 
	if(x==?20'b???10??1101?00???1?1) z |= 4'b0100; 
	if(x==?20'b?111?1??010??00??11?) z |= 4'b0100; 
	if(x==?20'b1???1??01?10??00?1?1) z |= 4'b1000; 
	if(x==?20'b??11?1??1011?00??11?) z |= 4'b0100; 
	if(x==?20'b????001?0?11?10?11??) z |= 4'b0100; 
	if(x==?20'b?11?0????111000???11) z |= 4'b0100; 
	if(x==?20'b???10??101?100???1?1) z |= 4'b0100; 
	if(x==?20'b1?1??1??1?11?0001??1) z |= 4'b1000; 
	if(x==?20'b?????10011?0?01?11??) z |= 4'b1000; 
	if(x==?20'b?????11??001??01110?) z |= 4'b1000; 
	if(x==?20'b?111???111??000?1??1) z |= 4'b0100; 
	if(x==?20'b?11?0?1??0??111???11) z |= 4'b0100; 
	if(x==?20'b11???1?1??10?101?1??) z |= 4'b1000; 
	if(x==?20'b111???1??010?00??11?) z |= 4'b1000; 
	if(x==?20'b???1???100??010??111) z |= 4'b0100; 
	if(x==?20'b11??1?0?100??0??11??) z |= 4'b1000; 
	if(x==?20'b?11101???10??00??11?) z |= 4'b0100; 
	if(x==?20'b1?1?1?0?100???0?11??) z |= 4'b1000; 
	if(x==?20'b???10?11111??0????01) z |= 4'b0100; 
	if(x==?20'b?11101??01???00??11?) z |= 4'b0100; 
	if(x==?20'b????001?0?11?01?11??) z |= 4'b0100; 
	if(x==?20'b111???10?01??00??11?) z |= 4'b1000; 
	if(x==?20'b1???1?????00?010?111) z |= 4'b1000; 
	if(x==?20'b1?1?1?101010?????1??) z |= 4'b1000; 
	if(x==?20'b????0011??1?010?11??) z |= 4'b0100; 
	if(x==?20'b?11??1?0??0??111??11) z |= 4'b1000; 
	if(x==?20'b111?1?????11?0001??1) z |= 4'b1000; 
	if(x==?20'b111???10??10?00??11?) z |= 4'b1000; 
	if(x==?20'b1???11?0?111??0???01) z |= 4'b1000; 
	if(x==?20'b?1?101?10101?????1??) z |= 4'b0100; 
	if(x==?20'b?1?1?0?1?001?0??11??) z |= 4'b0100; 
	if(x==?20'b1?1?1?111?0???0?1?11) z |= 4'b1000; 
	if(x==?20'b??1?011111??0?0?1?1?) z |= 4'b0100; 
	if(x==?20'b?1??011111??0?0?1?1?) z |= 4'b0100; 
	if(x==?20'b???10??101?1?10??11?) z |= 4'b0100; 
	if(x==?20'b????1100?1???01011??) z |= 4'b1000; 
	if(x==?20'b????111?111?111?????) z |= 4'b0010; 
	if(x==?20'b11?????1110???1?110?) z |= 4'b1000; 
	if(x==?20'b?1??0??100??01???111) z |= 4'b0100; 
	if(x==?20'b??111????011?1??110?) z |= 4'b0100; 
	if(x==?20'b?????1001?1??10011??) z |= 4'b1000; 
	if(x==?20'b?????11101?1?10?01??) z |= 4'b0100; 
	if(x==?20'b??1?0??100???11?1?11) z |= 4'b0100; 
	if(x==?20'b?111?1???10?000??11?) z |= 4'b0100; 
	if(x==?20'b?11???1?1101??00?11?) z |= 4'b1000; 
	if(x==?20'b?????0?1?00100??111?) z |= 4'b0100; 
	if(x==?20'b1???1??01?10?01??11?) z |= 4'b1000; 
	if(x==?20'b???1??11111?00????01) z |= 4'b0100; 
	if(x==?20'b??1?1110??11?0?01?1?) z |= 4'b1000; 
	if(x==?20'b?1??1110??11?0?01?1?) z |= 4'b1000; 
	if(x==?20'b?111?1??01??000??11?) z |= 4'b0100; 
	if(x==?20'b???10???0??1010??111) z |= 4'b0100; 
	if(x==?20'b?????1??1?00?1101?11) z |= 4'b1000; 
	if(x==?20'b?1?111?1?0?1?0??1?11) z |= 4'b0100; 
	if(x==?20'b???1??1?00??110?1?11) z |= 4'b0100; 
	if(x==?20'b?1??1?111110??0?1?1?) z |= 4'b1000; 
	if(x==?20'b??1?1??0??00??10?111) z |= 4'b1000; 
	if(x==?20'b111???1??01??000?11?) z |= 4'b1000; 
	if(x==?20'b?11??1??101100???11?) z |= 4'b0100; 
	if(x==?20'b????001??1?1001?11??) z |= 4'b0100; 
	if(x==?20'b1???1??01????101?111) z |= 4'b1000; 
	if(x==?20'b111???1???10?000?11?) z |= 4'b1000; 
	if(x==?20'b1???11???111??00??01) z |= 4'b1000; 
	if(x==?20'b1??????01??0?010?111) z |= 4'b1000; 
	if(x==?20'b??????1?00?1011?1?11) z |= 4'b0100; 
	if(x==?20'b????1?0?1?00??00111?) z |= 4'b1010; 
	if(x==?20'b??1?11?10111?0??1?1?) z |= 4'b0100; 
	if(x==?20'b1???1??0100??00?11??) z |= 4'b1000; 
	if(x==?20'b?????111?111?111????) z |= 4'b0001; 
	if(x==?20'b?1??1?????00?1101?11) z |= 4'b1000; 
	if(x==?20'b?11?1?0?100????011??) z |= 4'b1000; 
	if(x==?20'b??1?0?11111?0?????01) z |= 4'b0100; 
	if(x==?20'b??1????100??011?1?11) z |= 4'b0100; 
	if(x==?20'b???10??1???1101??111) z |= 4'b0100; 
	if(x==?20'b?1110?1?11?1??0?1??1) z |= 4'b0100; 
	if(x==?20'b?1??11?0?111???0??01) z |= 4'b1000; 
	if(x==?20'b???????0?100?100111?) z |= 4'b1000; 
	if(x==?20'b????11?01?10??1011??) z |= 4'b1000; 
	if(x==?20'b1?1?1?1011????10?1??) z |= 4'b1000; 
	if(x==?20'b??1???1?0101010??1??) z |= 4'b0100; 
	if(x==?20'b?11??0?1?0010???11??) z |= 4'b0100; 
	if(x==?20'b1????1????00?0111?11) z |= 4'b1000; 
	if(x==?20'b1?1??1111????000??11) z |= 4'b1000; 
	if(x==?20'b??1?0??101?101???11?) z |= 4'b0100; 
	if(x==?20'b?1??0??101?101???11?) z |= 4'b0100; 
	if(x==?20'b??1?1?11??0??0001?11) z |= 4'b1000; 
	if(x==?20'b111??1?01?11?0??1??1) z |= 4'b1000; 
	if(x==?20'b?11????11?01??00111?) z |= 4'b1000; 
	if(x==?20'b?1?101?1??1101???1??) z |= 4'b0100; 
	if(x==?20'b????0?110?110?1?11??) z |= 4'b0100; 
	if(x==?20'b??1?11?10???000?1?11) z |= 4'b0100; 
	if(x==?20'b?1??11?1?0??000?1?11) z |= 4'b0100; 
	if(x==?20'b?1?1111????1000???11) z |= 4'b0100; 
	if(x==?20'b?1??1???1?00??111?11) z |= 4'b1000; 
	if(x==?20'b?1??1?11???0?0001?11) z |= 4'b1000; 
	if(x==?20'b??1?1??01?10??10?11?) z |= 4'b1000; 
	if(x==?20'b?1??1??01?10??10?11?) z |= 4'b1000; 
	if(x==?20'b??1???111?0??0001?11) z |= 4'b1000; 
	if(x==?20'b?1????111?0??0001?11) z |= 4'b1000; 
	if(x==?20'b????1??01101??00?1?1) z |= 4'b1000; 
	if(x==?20'b?11??????011100?111?) z |= 4'b0100; 
	if(x==?20'b????0???001?001?111?) z |= 4'b0100; 
	if(x==?20'b???10??101??000??1?1) z |= 4'b0100; 
	if(x==?20'b?1???1??1010?010?1??) z |= 4'b1000; 
	if(x==?20'b?111??1?11?10?0?1??1) z |= 4'b0100; 
	if(x==?20'b1?1?11???11??0001?1?) z |= 4'b1000; 
	if(x==?20'b1???1??0??10?000?1?1) z |= 4'b1000; 
	if(x==?20'b?1?1??11?11?000?1?1?) z |= 4'b0100; 
	if(x==?20'b????0??1101100???1?1) z |= 4'b0100; 
	if(x==?20'b??1?11???0?1000?1?11) z |= 4'b0100; 
	if(x==?20'b?1??11???0?1000?1?11) z |= 4'b0100; 
	if(x==?20'b111??1??1?11?0?01??1) z |= 4'b1000; 
	if(x==?20'b111?1?10?1???1?1?1??) z |= 4'b1000; 
	if(x==?20'b????0?11010??10?11??) z |= 4'b0100; 
	if(x==?20'b?111101??1??01???1??) z |= 4'b0100; 
	if(x==?20'b111?1?0?100?????11??) z |= 4'b1000; 
	if(x==?20'b?11???10?101?00??11?) z |= 4'b1000; 
	if(x==?20'b?11?01??101??00??11?) z |= 4'b0100; 
	if(x==?20'b??110?11111???????01) z |= 4'b0100; 
	if(x==?20'b11?????1?10??10?110?) z |= 4'b1000; 
	if(x==?20'b??????101100?10?11??) z |= 4'b1000; 
	if(x==?20'b?????1?01?01?01011??) z |= 4'b1000; 
	if(x==?20'b11??11?0?111??????01) z |= 4'b1000; 
	if(x==?20'b?1?1?11?11?100??1?1?) z |= 4'b0100; 
	if(x==?20'b??11??1?0101?10??1??) z |= 4'b0100; 
	if(x==?20'b1???11??1100???01?1?) z |= 4'b1000; 
	if(x==?20'b?111?0?1?001????11??) z |= 4'b0100; 
	if(x==?20'b1?1?1?11??0??00?1?11) z |= 4'b1000; 
	if(x==?20'b?????11?100??01?110?) z |= 4'b0100; 
	if(x==?20'b1?1??11?1?11??001?1?) z |= 4'b1000; 
	if(x==?20'b??????11010?010?11??) z |= 4'b0100; 
	if(x==?20'b????11?0?010?01?11??) z |= 4'b1000; 
	if(x==?20'b?1?111?1?0???00?1?11) z |= 4'b0100; 
	if(x==?20'b????0?1101??010??11?) z |= 4'b0100; 
	if(x==?20'b1???1?1010?0??0?11??) z |= 4'b1000; 
	if(x==?20'b111??101??1???10?1??) z |= 4'b1000; 
	if(x==?20'b1???1??01101??0??1?1) z |= 4'b1000; 
	if(x==?20'b??11??11111?0?????01) z |= 4'b0100; 
	if(x==?20'b???101?10?01?0??11??) z |= 4'b0100; 
	if(x==?20'b????001??1?1100?11??) z |= 4'b0100; 
	if(x==?20'b???1??1100110???1?1?) z |= 4'b0100; 
	if(x==?20'b??111?1?01??010??1??) z |= 4'b0100; 
	if(x==?20'b11???1??1010?01??1??) z |= 4'b1000; 
	if(x==?20'b??????1?00?1110?1?11) z |= 4'b0100; 
	if(x==?20'b??1?1?????00?101?111) z |= 4'b1000; 
	if(x==?20'b11??11???111???0??01) z |= 4'b1000; 
	if(x==?20'b?1?????100??101??111) z |= 4'b0100; 
	if(x==?20'b???10?11111?00?????1) z |= 4'b0100; 
	if(x==?20'b???10??11011?0???1?1) z |= 4'b0100; 
	if(x==?20'b????01??0011?01?11??) z |= 4'b0100; 
	if(x==?20'b??????10110??10011??) z |= 4'b1000; 
	if(x==?20'b?1??11??0?1?000?1?11) z |= 4'b0100; 
	if(x==?20'b????0?110?1?010?11??) z |= 4'b0100; 
	if(x==?20'b??1???111110?00?1?1?) z |= 4'b1000; 
	if(x==?20'b1?1?110?101???0??1??) z |= 4'b1000; 
	if(x==?20'b?1????111110?00?1?1?) z |= 4'b1000; 
	if(x==?20'b?????1001?1??00111??) z |= 4'b1000; 
	if(x==?20'b?1?1?011?101?0???1??) z |= 4'b0100; 
	if(x==?20'b??1????100??110?1?11) z |= 4'b0100; 
	if(x==?20'b????11?0??10?010?11?) z |= 4'b1000; 
	if(x==?20'b????11???010?01011??) z |= 4'b1000; 
	if(x==?20'b??1?11??0111?00?1?1?) z |= 4'b0100; 
	if(x==?20'b?1??11??0111?00?1?1?) z |= 4'b0100; 
	if(x==?20'b??????1011?0?10011??) z |= 4'b1000; 
	if(x==?20'b?111???111?1?00?1??1) z |= 4'b0100; 
	if(x==?20'b1???11?0?111??00???1) z |= 4'b1000; 
	if(x==?20'b111?1???1?11?00?1??1) z |= 4'b1000; 
	if(x==?20'b?????1??1?00?0111?11) z |= 4'b1000; 
	if(x==?20'b1???1???1101??00?1?1) z |= 4'b1000; 
	if(x==?20'b11????101????101?1?1) z |= 4'b1000; 
	if(x==?20'b??111?11?1??101??1??) z |= 4'b0100; 
	if(x==?20'b?11?1???10??000?111?) z |= 4'b0100; 
	if(x==?20'b?11???110???111???11) z |= 4'b0100; 
	if(x==?20'b??1?0?1?111?00????01) z |= 4'b0100; 
	if(x==?20'b?1?101?1??1?010??1??) z |= 4'b0100; 
	if(x==?20'b?11???1?010101???1??) z |= 4'b0100; 
	if(x==?20'b????11?0??10?01011??) z |= 4'b1000; 
	if(x==?20'b1?1?1?10?1???010?1??) z |= 4'b1000; 
	if(x==?20'b?1?????1001?010?11??) z |= 4'b0100; 
	if(x==?20'b??110??1?001??0?11??) z |= 4'b0100; 
	if(x==?20'b11??11?1??1??101?1??) z |= 4'b1000; 
	if(x==?20'b????0?1??011010?11??) z |= 4'b0100; 
	if(x==?20'b??1????01??0?101?111) z |= 4'b1000; 
	if(x==?20'b11???1?1??10?010?1??) z |= 4'b1000; 
	if(x==?20'b???1???1101100???1?1) z |= 4'b0100; 
	if(x==?20'b??1?1????100?01011??) z |= 4'b1000; 
	if(x==?20'b?11????1??01?000111?) z |= 4'b1000; 
	if(x==?20'b??1101?????1101??1?1) z |= 4'b0100; 
	if(x==?20'b??1?011111?1??0?1?1?) z |= 4'b0100; 
	if(x==?20'b?1??0???0??1101??111) z |= 4'b0100; 
	if(x==?20'b?1??1?????00?0111?11) z |= 4'b1000; 
	if(x==?20'b?1???1?0?111??00??01) z |= 4'b1000; 
	if(x==?20'b?11?11?????0?111??11) z |= 4'b1000; 
	if(x==?20'b???101?1?0?10?0?11??) z |= 4'b0100; 
	if(x==?20'b????1??0?101?000?1?1) z |= 4'b1000; 
	if(x==?20'b111???1??101?00??11?) z |= 4'b1000; 
	if(x==?20'b?11???1??0?1111???11) z |= 4'b0100; 
	if(x==?20'b1?1??110?1???101?1??) z |= 4'b1000; 
	if(x==?20'b?11??1??1?0??111??11) z |= 4'b1000; 
	if(x==?20'b?111?1??101??00??11?) z |= 4'b0100; 
	if(x==?20'b???????01100??0011?1) z |= 4'b1000; 
	if(x==?20'b????0??1101?000??1?1) z |= 4'b0100; 
	if(x==?20'b????01??0?11001?11??) z |= 4'b0100; 
	if(x==?20'b????1??01?10?000?1?1) z |= 4'b1000; 
	if(x==?20'b111???1?1?10?00??11?) z |= 4'b1000; 
	if(x==?20'b1???1?101????01011??) z |= 4'b1000; 
	if(x==?20'b????01???011001?11??) z |= 4'b0100; 
	if(x==?20'b??110??101??0?0??1?1) z |= 4'b0100; 
	if(x==?20'b?11??1??1010??10?1??) z |= 4'b1000; 
	if(x==?20'b???101??00??00???111) z |= 4'b0100; 
	if(x==?20'b?111?1??01?1?00??11?) z |= 4'b0100; 
	if(x==?20'b1?????10??00??00?111) z |= 4'b1000; 
	if(x==?20'b????0??101?1000??1?1) z |= 4'b0100; 
	if(x==?20'b11??1??0??10?0?0?1?1) z |= 4'b1000; 
	if(x==?20'b??1?0??11?1?101??11?) z |= 4'b0100; 
	if(x==?20'b?1??0??11?1?101??11?) z |= 4'b0100; 
	if(x==?20'b??1?1??0?1?1?101?11?) z |= 4'b1000; 
	if(x==?20'b?1??1??0?1?1?101?11?) z |= 4'b1000; 
	if(x==?20'b????0???001100??11?1) z |= 4'b0100; 
	if(x==?20'b????0?11111??00???01) z |= 4'b0100; 
	if(x==?20'b??110011?1??0???1?1?) z |= 4'b0100; 
	if(x==?20'b??1110?1???1?10?11??) z |= 4'b0100; 
	if(x==?20'b??1?1?0?1?00?00?11??) z |= 4'b1000; 
	if(x==?20'b?1?111??0?1??00?1?11) z |= 4'b0100; 
	if(x==?20'b??1??11111?10?0?1?1?) z |= 4'b0100; 
	if(x==?20'b????0???001?100?111?) z |= 4'b0110; 
	if(x==?20'b?1??111?1?11?0?01?1?) z |= 4'b1000; 
	if(x==?20'b1???11?0??10?01??11?) z |= 4'b1000; 
	if(x==?20'b?1??1?0?10?0?00?11??) z |= 4'b1000; 
	if(x==?20'b111????11????0001?11) z |= 4'b1000; 
	if(x==?20'b???????01100?10?111?) z |= 4'b1000; 
	if(x==?20'b????11?0?111?00???01) z |= 4'b1000; 
	if(x==?20'b???1??11011?0?1?1?1?) z |= 4'b0100; 
	if(x==?20'b1???1??01????010?111) z |= 4'b1000; 
	if(x==?20'b???10??1???1010??111) z |= 4'b0100; 
	if(x==?20'b??1????100?1?11?1?11) z |= 4'b0100; 
	if(x==?20'b???????0?100?001111?) z |= 4'b1001; 
	if(x==?20'b??1?1?111?0??00?1?11) z |= 4'b1000; 
	if(x==?20'b???10??1??110?1?1?11) z |= 4'b0100; 
	if(x==?20'b?1???0?1?001?00?11??) z |= 4'b0100; 
	if(x==?20'b??110?1?111??0????01) z |= 4'b0100; 
	if(x==?20'b1?1????0?100?1??111?) z |= 4'b1000; 
	if(x==?20'b?111?1??00??01???1?1) z |= 4'b0100; 
	if(x==?20'b?1??1?111??0?00?1?11) z |= 4'b1000; 
	if(x==?20'b?1?10???001??1??111?) z |= 4'b0100; 
	if(x==?20'b1?1?1?11?11??00?1?1?) z |= 4'b1000; 
	if(x==?20'b??????11111?000???01) z |= 4'b0100; 
	if(x==?20'b?1?111?1?11??00?1?1?) z |= 4'b0100; 
	if(x==?20'b?1??0?1101??01???11?) z |= 4'b0100; 
	if(x==?20'b??1?11?10??1?00?1?11) z |= 4'b0100; 
	if(x==?20'b?1??11?1?0?1?00?1?11) z |= 4'b0100; 
	if(x==?20'b11???1?0?111??0???01) z |= 4'b1000; 
	if(x==?20'b1?1????0?100??1?111?) z |= 4'b1000; 
	if(x==?20'b111???1???00??10?1?1) z |= 4'b1000; 
	if(x==?20'b1???1??0?101?00??1?1) z |= 4'b1000; 
	if(x==?20'b?1????1?00??011?1?11) z |= 4'b0100; 
	if(x==?20'b????????1100?100111?) z |= 4'b1000; 
	if(x==?20'b????11???111?000??01) z |= 4'b1000; 
	if(x==?20'b1???1??01?10?00??1?1) z |= 4'b1000; 
	if(x==?20'b???10??1101??00??1?1) z |= 4'b0100; 
	if(x==?20'b??1??1????00?1101?11) z |= 4'b1000; 
	if(x==?20'b?1?10???001???1?111?) z |= 4'b0100; 
	if(x==?20'b????0???0011?01?111?) z |= 4'b0100; 
	if(x==?20'b???10??101?1?00??1?1) z |= 4'b0100; 
	if(x==?20'b??1???11?101010??1??) z |= 4'b0100; 
	if(x==?20'b??11??1?111?00????01) z |= 4'b0100; 
	if(x==?20'b???????0110??100111?) z |= 4'b1000; 
	if(x==?20'b?1???1?0??0??1101?11) z |= 4'b1000; 
	if(x==?20'b??110?11111?0??????1) z |= 4'b0100; 
	if(x==?20'b??1?0?1??0??011?1?11) z |= 4'b0100; 
	if(x==?20'b1???1???10?0?0?0111?) z |= 4'b1000; 
	if(x==?20'b???10?1?011?00??1??1) z |= 4'b0100; 
	if(x==?20'b???????011?0?100111?) z |= 4'b1000; 
	if(x==?20'b?1?1?11111?1?0??1?1?) z |= 4'b0100; 
	if(x==?20'b?1??11??101??010?1??) z |= 4'b1000; 
	if(x==?20'b1???11??11?0?0?11?1?) z |= 4'b1000; 
	if(x==?20'b1?1?1?101??0???0?11?) z |= 4'b1000; 
	if(x==?20'b1?1?111?1?11??0?1?1?) z |= 4'b1000; 
	if(x==?20'b???1??110?111?0?1?1?) z |= 4'b0100; 
	if(x==?20'b11??11?0?111???0???1) z |= 4'b1000; 
	if(x==?20'b11???1???111??00??01) z |= 4'b1000; 
	if(x==?20'b???1???10?010?0?111?) z |= 4'b0100; 
	if(x==?20'b1????1?0?110??001??1) z |= 4'b1000; 
	if(x==?20'b1???1????101?000?1?1) z |= 4'b1000; 
	if(x==?20'b1???1???1?10?000?1?1) z |= 4'b1000; 
	if(x==?20'b???1???1101?000??1?1) z |= 4'b0100; 
	if(x==?20'b??11?10????1001?11??) z |= 4'b0100; 
	if(x==?20'b????????0011001?111?) z |= 4'b0100; 
	if(x==?20'b?1?101?10??10????11?) z |= 4'b0100; 
	if(x==?20'b???1???101?1000??1?1) z |= 4'b0100; 
	if(x==?20'b111?1?1?11???1?1?1??) z |= 4'b1000; 
	if(x==?20'b?1??0??100???10??111) z |= 4'b0100; 
	if(x==?20'b??????10110??00111??) z |= 4'b1000; 
	if(x==?20'b??11011?00??0???1?1?) z |= 4'b0100; 
	if(x==?20'b?11?1????01?10??110?) z |= 4'b0100; 
	if(x==?20'b?11???1?1101?00??11?) z |= 4'b1000; 
	if(x==?20'b11???110??00???01?1?) z |= 4'b1000; 
	if(x==?20'b????11?01??1?10011??) z |= 4'b1000; 
	if(x==?20'b???1??11111??00???01) z |= 4'b0100; 
	if(x==?20'b????0???0?11001?111?) z |= 4'b0100; 
	if(x==?20'b????0????011001?111?) z |= 4'b0100; 
	if(x==?20'b?11?1?1?01??101??1??) z |= 4'b0100; 
	if(x==?20'b??????1011?0?00111??) z |= 4'b1000; 
	if(x==?20'b????01??0?11100?11??) z |= 4'b0100; 
	if(x==?20'b??1?1??0??00?01??111) z |= 4'b1000; 
	if(x==?20'b????01???011100?11??) z |= 4'b0100; 
	if(x==?20'b?11????1?10???01110?) z |= 4'b1000; 
	if(x==?20'b??1?1??0?101??00?1?1) z |= 4'b1000; 
	if(x==?20'b???1011101??0????11?) z |= 4'b0100; 
	if(x==?20'b?1??0??1101?00???1?1) z |= 4'b0100; 
	if(x==?20'b???????0?100?00011?1) z |= 4'b1000; 
	if(x==?20'b??1?1??01?10??00?1?1) z |= 4'b1000; 
	if(x==?20'b1???11???111?00???01) z |= 4'b1000; 
	if(x==?20'b????1110?0?1??0111??) z |= 4'b1000; 
	if(x==?20'b?1110??101??0????1?1) z |= 4'b0100; 
	if(x==?20'b?11??1??1011?00??11?) z |= 4'b0100; 
	if(x==?20'b?1??0??101?100???1?1) z |= 4'b0100; 
	if(x==?20'b????0???001?000?11?1) z |= 4'b0100; 
	if(x==?20'b1???1110??10???0?11?) z |= 4'b1000; 
	if(x==?20'b111?1??0??10???0?1?1) z |= 4'b1000; 
	if(x==?20'b?11??1?1??10?101?1??) z |= 4'b1000; 
	if(x==?20'b??110???01??000??1?1) z |= 4'b0100; 
	if(x==?20'b?1?????100??010??111) z |= 4'b0100; 
	if(x==?20'b??11???11011?1???11?) z |= 4'b0100; 
	if(x==?20'b1???1??011???0?11?11) z |= 4'b1000; 
	if(x==?20'b11??1???1101??1??11?) z |= 4'b1000; 
	if(x==?20'b?1??0?11111??0????01) z |= 4'b0100; 
	if(x==?20'b??1?0?11111???0???01) z |= 4'b0100; 
	if(x==?20'b??1111????1111??1??1) z |= 4'b0100; 
	if(x==?20'b????0?110?11?10?11??) z |= 4'b0100; 
	if(x==?20'b??1?1?????00?010?111) z |= 4'b1000; 
	if(x==?20'b11?????0??10?000?1?1) z |= 4'b1000; 
	if(x==?20'b??1?0?1?011??11?1?1?) z |= 4'b0100; 
	if(x==?20'b?1??11?0?111?0????01) z |= 4'b1000; 
	if(x==?20'b????11?01?10?01?11??) z |= 4'b1000; 
	if(x==?20'b1?1?1?1011???01??1??) z |= 4'b1000; 
	if(x==?20'b??1?11?0?111??0???01) z |= 4'b1000; 
	if(x==?20'b??111?11?1??010??1??) z |= 4'b0100; 
	if(x==?20'b?1???1?0?110?11?1?1?) z |= 4'b1000; 
	if(x==?20'b??1?0??101?1?10??11?) z |= 4'b0100; 
	if(x==?20'b?1??0??101?1?10??11?) z |= 4'b0100; 
	if(x==?20'b?11????11?01?00?111?) z |= 4'b1000; 
	if(x==?20'b?1?1?01??0??000??11?) z |= 4'b0100; 
	if(x==?20'b?11????1110???1?110?) z |= 4'b1000; 
	if(x==?20'b11????1111????111??1) z |= 4'b1000; 
	if(x==?20'b?11?1????011?1??110?) z |= 4'b0100; 
	if(x==?20'b?1?101?1??11?10??1??) z |= 4'b0100; 
	if(x==?20'b1????11011?0???01?1?) z |= 4'b1000; 
	if(x==?20'b1???11???110?0?11?1?) z |= 4'b1000; 
	if(x==?20'b?????11??010?10011??) z |= 4'b1000; 
	if(x==?20'b?????11?010?001?11??) z |= 4'b0100; 
	if(x==?20'b??1?1??01?10?01??11?) z |= 4'b1000; 
	if(x==?20'b?1??1??01?10?01??11?) z |= 4'b1000; 
	if(x==?20'b????1??01101?00??1?1) z |= 4'b1000; 
	if(x==?20'b??1101?????1010??1?1) z |= 4'b0100; 
	if(x==?20'b?1????11111?00????01) z |= 4'b0100; 
	if(x==?20'b??1???11111?0?0???01) z |= 4'b0100; 
	if(x==?20'b11????101????010?1?1) z |= 4'b1000; 
	if(x==?20'b?1??0???0??1010??111) z |= 4'b0100; 
	if(x==?20'b?1????1?00??110?1?11) z |= 4'b0100; 
	if(x==?20'b??????110?11010?11??) z |= 4'b0100; 
	if(x==?20'b???1011?0?110???1?1?) z |= 4'b0100; 
	if(x==?20'b?1??11???111?0?0??01) z |= 4'b1000; 
	if(x==?20'b??1?1??01????101?111) z |= 4'b1000; 
	if(x==?20'b?1110??10???00????11) z |= 4'b0100; 
	if(x==?20'b????11??1?10?01011??) z |= 4'b1000; 
	if(x==?20'b1?1?1?1?11???010?1??) z |= 4'b1000; 
	if(x==?20'b11??11?1??1??010?1??) z |= 4'b1000; 
	if(x==?20'b??1?11???111??00??01) z |= 4'b1000; 
	if(x==?20'b??1????01??0?010?111) z |= 4'b1000; 
	if(x==?20'b111?1??0???0??00??11) z |= 4'b1000; 
	if(x==?20'b????0?11111?000????1) z |= 4'b0100; 
	if(x==?20'b????0??11011?00??1?1) z |= 4'b0100; 
	if(x==?20'b??1?0?1??0??110?1?11) z |= 4'b0100; 
	if(x==?20'b??1????1010100??11??) z |= 4'b0100; 
	if(x==?20'b?1??1???1010??0011??) z |= 4'b1000; 
	if(x==?20'b??1?1??0100??00?11??) z |= 4'b1000; 
	if(x==?20'b???1101??1??000??11?) z |= 4'b0100; 
	if(x==?20'b??11??1111??11??1?1?) z |= 4'b0100; 
	if(x==?20'b?1?1?1?1??11010??1??) z |= 4'b0100; 
	if(x==?20'b??1?0?1??11?011?1?1?) z |= 4'b0100; 
	if(x==?20'b?111101??1???10??1??) z |= 4'b0100; 
	if(x==?20'b????11?0?111?000???1) z |= 4'b1000; 
	if(x==?20'b?1???1?0?11??1101?1?) z |= 4'b1000; 
	if(x==?20'b?????1?01110??001??1) z |= 4'b1000; 
	if(x==?20'b?1??0??1???1101??111) z |= 4'b0100; 
	if(x==?20'b????1???1101?000?1?1) z |= 4'b1000; 
	if(x==?20'b????0?1?011100??1??1) z |= 4'b0100; 
	if(x==?20'b1?1?1?10???0?0?0?11?) z |= 4'b1000; 
	if(x==?20'b??110?1?111?00?????1) z |= 4'b0100; 
	if(x==?20'b?1?101?10???0?0??11?) z |= 4'b0100; 
	if(x==?20'b????0?11??11001?11??) z |= 4'b0100; 
	if(x==?20'b1????101??1??000?11?) z |= 4'b1000; 
	if(x==?20'b????????1100?001111?) z |= 4'b1000; 
	if(x==?20'b11???01?1????00111??) z |= 4'b1000; 
	if(x==?20'b??1??1????00?0111?11) z |= 4'b1000; 
	if(x==?20'b????????0011100?111?) z |= 4'b0100; 
	if(x==?20'b?1?1?11?11?1?00?1?1?) z |= 4'b0100; 
	if(x==?20'b1???11??1100??0?1?1?) z |= 4'b1000; 
	if(x==?20'b??1?0??1011?00??1??1) z |= 4'b0100; 
	if(x==?20'b???????11011000??1?1) z |= 4'b0100; 
	if(x==?20'b???????0110??001111?) z |= 4'b1000; 
	if(x==?20'b1?1??11?1?11?00?1?1?) z |= 4'b1000; 
	if(x==?20'b?1??1??0?110??001??1) z |= 4'b1000; 
	if(x==?20'b?1???1?0??0??0111?11) z |= 4'b1000; 
	if(x==?20'b11???1?0?111??00???1) z |= 4'b1000; 
	if(x==?20'b???11?1101??0?0??11?) z |= 4'b0100; 
	if(x==?20'b????0???0?11100?111?) z |= 4'b0100; 
	if(x==?20'b??111??1???1010?11??) z |= 4'b0100; 
	if(x==?20'b????0????011100?111?) z |= 4'b0100; 
	if(x==?20'b???????011?0?001111?) z |= 4'b1000; 
	if(x==?20'b111??101??1??01??1??) z |= 4'b1000; 
	if(x==?20'b?1?1??11111??0????01) z |= 4'b0100; 
	if(x==?20'b11??1??11????01011??) z |= 4'b1000; 
	if(x==?20'b??1?0?1?11??00??1?01) z |= 4'b0100; 
	if(x==?20'b??11??11111???0???01) z |= 4'b0100; 
	if(x==?20'b???1?1??0?110?1?1?11) z |= 4'b0100; 
	if(x==?20'b?1??0??101??000??1?1) z |= 4'b0100; 
	if(x==?20'b??????10??00?000?111) z |= 4'b1000; 
	if(x==?20'b????01??00??000??111) z |= 4'b0100; 
	if(x==?20'b1???11?1??10?0?0?11?) z |= 4'b1000; 
	if(x==?20'b???1??110011?0??1?1?) z |= 4'b0100; 
	if(x==?20'b??1101??1???010?11??) z |= 4'b0100; 
	if(x==?20'b11??11???111?0????01) z |= 4'b1000; 
	if(x==?20'b??1?1??0??10?000?1?1) z |= 4'b1000; 
	if(x==?20'b1?1?11???111??0???01) z |= 4'b1000; 
	if(x==?20'b11??11????11??111?1?) z |= 4'b1000; 
	if(x==?20'b???10?11111??00????1) z |= 4'b0100; 
	if(x==?20'b?1110???01??00???1?1) z |= 4'b0100; 
	if(x==?20'b??111???0???010?11?1) z |= 4'b0100; 
	if(x==?20'b????11?01??1?00111??) z |= 4'b1000; 
	if(x==?20'b?1???1?0??11??001?01) z |= 4'b1000; 
	if(x==?20'b1???11??110???001?1?) z |= 4'b1000; 
	if(x==?20'b1???11?0?111?00????1) z |= 4'b1000; 
	if(x==?20'b?11?0?11111???????01) z |= 4'b0100; 
	if(x==?20'b11??????1100??1?111?) z |= 4'b1000; 
	if(x==?20'b?11????1?10??10?110?) z |= 4'b1000; 
	if(x==?20'b1????1?01110??0?1??1) z |= 4'b1000; 
	if(x==?20'b??11????0011?1??111?) z |= 4'b0100; 
	if(x==?20'b1???1???1101?00??1?1) z |= 4'b1000; 
	if(x==?20'b???10?1?0111?0??1??1) z |= 4'b0100; 
	if(x==?20'b1?1????1???0?10011?1) z |= 4'b1000; 
	if(x==?20'b111????0??10??00?1?1) z |= 4'b1000; 
	if(x==?20'b?11?11?0?111??????01) z |= 4'b1000; 
	if(x==?20'b??1?0?1?111??00???01) z |= 4'b0100; 
	if(x==?20'b11????10???1?01011??) z |= 4'b1000; 
	if(x==?20'b?1?11???0???001?11?1) z |= 4'b0100; 
	if(x==?20'b?1?101?????1001?11??) z |= 4'b0100; 
	if(x==?20'b?11???1?0101?10??1??) z |= 4'b0100; 
	if(x==?20'b??1?11??1100???01?1?) z |= 4'b1000; 
	if(x==?20'b???10110????000?1??1) z |= 4'b0100; 
	if(x==?20'b?1???1??1?0??1101?11) z |= 4'b1000; 
	if(x==?20'b?????11?010?100?11??) z |= 4'b0100; 
	if(x==?20'b11???1101?00????1?1?) z |= 4'b1000; 
	if(x==?20'b???1??11111?000????1) z |= 4'b0100; 
	if(x==?20'b???1???11011?00??1?1) z |= 4'b0100; 
	if(x==?20'b11?????1???0?01011?1) z |= 4'b1000; 
	if(x==?20'b???1??11?01100??1?1?) z |= 4'b0100; 
	if(x==?20'b??110?????110?1?1?11) z |= 4'b0100; 
	if(x==?20'b?1???1?0?111?00???01) z |= 4'b1000; 
	if(x==?20'b?11?1????01??01?110?) z |= 4'b0100; 
	if(x==?20'b1????1?0111???00??11) z |= 4'b1000; 
	if(x==?20'b?11101?????101???1?1) z |= 4'b0100; 
	if(x==?20'b??1?1??01101??0??1?1) z |= 4'b1000; 
	if(x==?20'b1???11???111?000???1) z |= 4'b1000; 
	if(x==?20'b?11???11111?0?????01) z |= 4'b0100; 
	if(x==?20'b??11011?00?1????1?1?) z |= 4'b0100; 
	if(x==?20'b???????01100?00?11?1) z |= 4'b1000; 
	if(x==?20'b??1???1??0?1011?1?11) z |= 4'b0100; 
	if(x==?20'b111???101?????10?1?1) z |= 4'b1000; 
	if(x==?20'b1????1??1110??001??1) z |= 4'b1000; 
	if(x==?20'b???10?1??11100????11) z |= 4'b0100; 
	if(x==?20'b?11??1??1010?01??1??) z |= 4'b1000; 
	if(x==?20'b?1????1100110???1?1?) z |= 4'b0100; 
	if(x==?20'b?11?1?1?01??010??1??) z |= 4'b0100; 
	if(x==?20'b???1??1?011100??1??1) z |= 4'b0100; 
	if(x==?20'b1?????10??00?00??111) z |= 4'b1000; 
	if(x==?20'b?111????00??000???11) z |= 4'b0100; 
	if(x==?20'b111???????00?000??11) z |= 4'b1000; 
	if(x==?20'b???101??00???00??111) z |= 4'b0100; 
	if(x==?20'b?11?11???111???0??01) z |= 4'b1000; 
	if(x==?20'b??1???1?111?000???01) z |= 4'b0100; 
	if(x==?20'b?1???????100?100111?) z |= 4'b1000; 
	if(x==?20'b11????1111???11?1??1) z |= 4'b1000; 
	if(x==?20'b111?11?1??1???10?1??) z |= 4'b1000; 
	if(x==?20'b?1??0?11111?00?????1) z |= 4'b0100; 
	if(x==?20'b?1??0??11011?0???1?1) z |= 4'b0100; 
	if(x==?20'b??1?0?11111?0?0????1) z |= 4'b0100; 
	if(x==?20'b??????1100??111???11) z |= 4'b0100; 
	if(x==?20'b1????1111?0??0?0??11) z |= 4'b1000; 
	if(x==?20'b??1?0?1??11?110?1?1?) z |= 4'b0100; 
	if(x==?20'b11???11?1?00???01?1?) z |= 4'b1000; 
	if(x==?20'b?11?1??0100??0??11??) z |= 4'b1000; 
	if(x==?20'b??110011?1???0??1?1?) z |= 4'b0100; 
	if(x==?20'b????0?1?011?000?1??1) z |= 4'b0100; 
	if(x==?20'b????0???0011?00?11?1) z |= 4'b0100; 
	if(x==?20'b?????11??010?00111??) z |= 4'b1000; 
	if(x==?20'b??110011?1????0?1?1?) z |= 4'b0100; 
	if(x==?20'b?1??11?0?111?0?0???1) z |= 4'b1000; 
	if(x==?20'b?1???1???111?000??01) z |= 4'b1000; 
	if(x==?20'b11??1100??1??0??1?1?) z |= 4'b1000; 
	if(x==?20'b??1?11?0?111??00???1) z |= 4'b1000; 
	if(x==?20'b?1???1?01110???01??1) z |= 4'b1000; 
	if(x==?20'b1????1111??0??00??11) z |= 4'b1000; 
	if(x==?20'b11??1100??1???0?1?1?) z |= 4'b1000; 
	if(x==?20'b?????1?0?110?0001??1) z |= 4'b1000; 
	if(x==?20'b????11?100??00??1?11) z |= 4'b0100; 
	if(x==?20'b???1111?0??100????11) z |= 4'b0100; 
	if(x==?20'b????1?11??00??001?11) z |= 4'b1000; 
	if(x==?20'b??1?1???1101??00?1?1) z |= 4'b1000; 
	if(x==?20'b??1111????11?11?1??1) z |= 4'b0100; 
	if(x==?20'b?11???101????101?1?1) z |= 4'b1000; 
	if(x==?20'b????11????00?111??11) z |= 4'b1000; 
	if(x==?20'b????0?11??11100?11??) z |= 4'b0100; 
	if(x==?20'b1???1??011????001?11) z |= 4'b1000; 
	if(x==?20'b??11?11?00?10???1?1?) z |= 4'b0100; 
	if(x==?20'b???1111??0?10?0???11) z |= 4'b0100; 
	if(x==?20'b????????1100?00011?1) z |= 4'b1000; 
	if(x==?20'b?11?1?11?1??101??1??) z |= 4'b0100; 
	if(x==?20'b??1?0?1?01110???1??1) z |= 4'b0100; 
	if(x==?20'b??1?????001?001?111?) z |= 4'b0100; 
	if(x==?20'b1?????1???00?000?111) z |= 4'b1000; 
	if(x==?20'b???1?1??00??000??111) z |= 4'b0100; 
	if(x==?20'b?11?0??1?001??0?11??) z |= 4'b0100; 
	if(x==?20'b?11?11?1??1??101?1??) z |= 4'b1000; 
	if(x==?20'b1?1??1?0??0??000?11?) z |= 4'b1000; 
	if(x==?20'b?11??1?1??10?010?1??) z |= 4'b1000; 
	if(x==?20'b?111?1??00???10??1?1) z |= 4'b0100; 
	if(x==?20'b??????111?00??001?11) z |= 4'b1000; 
	if(x==?20'b?1?????1101100???1?1) z |= 4'b0100; 
	if(x==?20'b?11?01?????1101??1?1) z |= 4'b0100; 
	if(x==?20'b????0111?10??01?11??) z |= 4'b0100; 
	if(x==?20'b????11??00?100??1?11) z |= 4'b0100; 
	if(x==?20'b????????0011000?11?1) z |= 4'b0100; 
	if(x==?20'b1?????1?11?0?0?11?11) z |= 4'b1000; 
	if(x==?20'b?1???1?0?11??0111?1?) z |= 4'b1000; 
	if(x==?20'b1???11???110??001?1?) z |= 4'b1000; 
	if(x==?20'b111???1???00?01??1?1) z |= 4'b1000; 
	if(x==?20'b?1??1?101????01011??) z |= 4'b1000; 
	if(x==?20'b?11?0??101??0?0??1?1) z |= 4'b0100; 
	if(x==?20'b??1?01?1???1010?11??) z |= 4'b0100; 
	if(x==?20'b?1??01??00??00???111) z |= 4'b0100; 
	if(x==?20'b??1???10??00??00?111) z |= 4'b1000; 
	if(x==?20'b?11?1??0??10?0?0?1?1) z |= 4'b1000; 
	if(x==?20'b????111??01??10011??) z |= 4'b1000; 
	if(x==?20'b11???????100?10?111?) z |= 4'b1000; 
	if(x==?20'b??1?111?111??00???10) z |= 4'b1100; 
	if(x==?20'b??11??1?111??00???01) z |= 4'b0100; 
	if(x==?20'b11???110110??0??1???) z |= 4'b1000; 
	if(x==?20'b?1?10?11111??0?????1) z |= 4'b0100; 
	if(x==?20'b11???110110???0?1???) z |= 4'b1000; 
	if(x==?20'b??110?11111???0????1) z |= 4'b0100; 
	if(x==?20'b1?1??101?????000?11?) z |= 4'b1000; 
	if(x==?20'b?11?0011?1??0???1?1?) z |= 4'b0100; 
	if(x==?20'b??11??1111???11?1?1?) z |= 4'b0100; 
	if(x==?20'b?????111?10?001?11??) z |= 4'b0100; 
	if(x==?20'b???10?1?011??00?1??1) z |= 4'b0100; 
	if(x==?20'b1?1?1?101??0?0???11?) z |= 4'b1000; 
	if(x==?20'b?11?1100???0?0??1?1?) z |= 4'b1000; 
	if(x==?20'b?11?1100??1????01?1?) z |= 4'b1000; 
	if(x==?20'b1?1?11??110????01?1?) z |= 4'b1000; 
	if(x==?20'b1?????1??101?000?11?) z |= 4'b1000; 
	if(x==?20'b11??11?0?111?0?????1) z |= 4'b1000; 
	if(x==?20'b?1????1101??010??11?) z |= 4'b0100; 
	if(x==?20'b???1?1??101?000??11?) z |= 4'b0100; 
	if(x==?20'b11???1???111?00???01) z |= 4'b1000; 
	if(x==?20'b1?1?11?0?111??0????1) z |= 4'b1000; 
	if(x==?20'b????11?0111??0?0??11) z |= 4'b1000; 
	if(x==?20'b111???1???00?0?0??11) z |= 4'b1000; 
	if(x==?20'b11?????011???0001??1) z |= 4'b1000; 
	if(x==?20'b1?????1?1?10?000?11?) z |= 4'b1000; 
	if(x==?20'b?1????11011?0?1?1?1?) z |= 4'b0100; 
	if(x==?20'b??1?1??01????010?111) z |= 4'b1000; 
	if(x==?20'b1????1?0?110?00?1??1) z |= 4'b1000; 
	if(x==?20'b?1??0??1???1010??111) z |= 4'b0100; 
	if(x==?20'b?1???111?111?00???10) z |= 4'b1100; 
	if(x==?20'b1???1?11??00??0?1?11) z |= 4'b1000; 
	if(x==?20'b???111?100???0??1?11) z |= 4'b0100; 
	if(x==?20'b?????11?110??01011??) z |= 4'b1000; 
	if(x==?20'b?111?1??00??0?0???11) z |= 4'b0100; 
	if(x==?20'b????1???001?000?111?) z |= 4'b0100; 
	if(x==?20'b???1?1??01?1000??11?) z |= 4'b0100; 
	if(x==?20'b?1??0??1??110?1?1?11) z |= 4'b0100; 
	if(x==?20'b?1?11???0???100?11?1) z |= 4'b0100; 
	if(x==?20'b111?1???1??0??00??11) z |= 4'b1000; 
	if(x==?20'b??11????001??01?111?) z |= 4'b0100; 
	if(x==?20'b1?1???101????00111??) z |= 4'b1000; 
	if(x==?20'b?11?0?1?111??0????01) z |= 4'b0100; 
	if(x==?20'b11??11????11?11?1?1?) z |= 4'b1000; 
	if(x==?20'b?11?01111110????1???) z |= 4'b1100; 
	if(x==?20'b?????11??011010?11??) z |= 4'b0100; 
	if(x==?20'b?1??1??01110??0?1??1) z |= 4'b1000; 
	if(x==?20'b??11011??011?0??1???) z |= 4'b0100; 
	if(x==?20'b??11????00??000?1?11) z |= 4'b0100; 
	if(x==?20'b?1?101?10??1??0??11?) z |= 4'b0100; 
	if(x==?20'b11????????00?0001?11) z |= 4'b1000; 
	if(x==?20'b?1111???0???0?1?11?1) z |= 4'b0100; 
	if(x==?20'b?11?11100111????1???) z |= 4'b1100; 
	if(x==?20'b11?????011???0?11?11) z |= 4'b1000; 
	if(x==?20'b??11011??011??0?1???) z |= 4'b0100; 
	if(x==?20'b??11?1???0?10?1?1?11) z |= 4'b0100; 
	if(x==?20'b1?????111?00??0?1?11) z |= 4'b1000; 
	if(x==?20'b????0?11?1110?0???11) z |= 4'b0100; 
	if(x==?20'b?111???10??100????11) z |= 4'b0100; 
	if(x==?20'b111?1??01?????00??11) z |= 4'b1000; 
	if(x==?20'b??11011?00???0??1?1?) z |= 4'b0100; 
	if(x==?20'b?1?1??11111?00?????1) z |= 4'b0100; 
	if(x==?20'b11???110??00?0??1?1?) z |= 4'b1000; 
	if(x==?20'b??110?????11000?1??1) z |= 4'b0100; 
	if(x==?20'b??11??11111?0?0????1) z |= 4'b0100; 
	if(x==?20'b??11011?00????0?1?1?) z |= 4'b0100; 
	if(x==?20'b111?1??0111???0????1) z |= 4'b1000; 
	if(x==?20'b11???110??00??0?1?1?) z |= 4'b1000; 
	if(x==?20'b??1?0??10111?0??1??1) z |= 4'b0100; 
	if(x==?20'b111????1???0??1011?1) z |= 4'b1000; 
	if(x==?20'b???1??1?011?000?1??1) z |= 4'b0100; 
	if(x==?20'b???111??00?1?0??1?11) z |= 4'b0100; 
	if(x==?20'b??1?11????10?010?11?) z |= 4'b1000; 
	if(x==?20'b1?1?1?1?1??0?0?0?11?) z |= 4'b1000; 
	if(x==?20'b?11??1?0?111??0???01) z |= 4'b1000; 
	if(x==?20'b??1???1??0?1110?1?11) z |= 4'b0100; 
	if(x==?20'b???????1?100?000111?) z |= 4'b1001; 
	if(x==?20'b11??11???111?0?0???1) z |= 4'b1000; 
	if(x==?20'b??1?1??0?101?00??1?1) z |= 4'b1000; 
	if(x==?20'b1?1?11???111??00???1) z |= 4'b1000; 
	if(x==?20'b???1011101????0??11?) z |= 4'b0100; 
	if(x==?20'b??1?1??01?10?00??1?1) z |= 4'b1000; 
	if(x==?20'b1????1???110?0001??1) z |= 4'b1000; 
	if(x==?20'b1?1????1???0?00111?1) z |= 4'b1000; 
	if(x==?20'b?1110??1???100????11) z |= 4'b0100; 
	if(x==?20'b?1??0??1101??00??1?1) z |= 4'b0100; 
	if(x==?20'b111???1?1????101?1?1) z |= 4'b1000; 
	if(x==?20'b?1????101?00?00?11??) z |= 4'b1000; 
	if(x==?20'b?1??1??0111???00??11) z |= 4'b1000; 
	if(x==?20'b?1110??101????0??1?1) z |= 4'b0100; 
	if(x==?20'b1?1?1?101????0?0?11?) z |= 4'b1000; 
	if(x==?20'b?1110??1?111?0?????1) z |= 4'b0100; 
	if(x==?20'b?1??0??101?1?00??1?1) z |= 4'b0100; 
	if(x==?20'b?11???1?111?00????01) z |= 4'b0100; 
	if(x==?20'b111?1??0??10?0???1?1) z |= 4'b1000; 
	if(x==?20'b?1??1???1110??001??1) z |= 4'b1000; 
	if(x==?20'b?1?1?1?10??10?0??11?) z |= 4'b0100; 
	if(x==?20'b?1???1??1?0??0111?11) z |= 4'b1000; 
	if(x==?20'b?11?0?11111?0??????1) z |= 4'b0100; 
	if(x==?20'b??1?01???001?00?11??) z |= 4'b0100; 
	if(x==?20'b1?1??1111?0????0??11) z |= 4'b1000; 
	if(x==?20'b??1?1???10?0?0?0111?) z |= 4'b1000; 
	if(x==?20'b1???111?111???00??1?) z |= 4'b1000; 
	if(x==?20'b???1111?0???000???11) z |= 4'b0100; 
	if(x==?20'b?1??0?1?011?00??1??1) z |= 4'b0100; 
	if(x==?20'b?111?1?????1101??1?1) z |= 4'b0100; 
	if(x==?20'b?1?1??11??110?1?1?1?) z |= 4'b0100; 
	if(x==?20'b??1?0?1?011?0?0?1??1) z |= 4'b0100; 
	if(x==?20'b??1?0??1?11100????11) z |= 4'b0100; 
	if(x==?20'b111?1???111???00???1) z |= 4'b1000; 
	if(x==?20'b??1?11??11?0?0?11?1?) z |= 4'b1000; 
	if(x==?20'b??1????1011100??1??1) z |= 4'b0100; 
	if(x==?20'b??1?0?1?111?000????1) z |= 4'b0100; 
	if(x==?20'b?11?11?0?111???0???1) z |= 4'b1000; 
	if(x==?20'b?1????110?111?0?1?1?) z |= 4'b0100; 
	if(x==?20'b?11??1???111??00??01) z |= 4'b1000; 
	if(x==?20'b11???1111??0???0??11) z |= 4'b1000; 
	if(x==?20'b?1???1?0?110?0?01??1) z |= 4'b1000; 
	if(x==?20'b?1??1?11??00???01?11) z |= 4'b1000; 
	if(x==?20'b1????111???0?000??11) z |= 4'b1000; 
	if(x==?20'b?1?????10?010?0?111?) z |= 4'b0100; 
	if(x==?20'b?1?101?1???10?0??11?) z |= 4'b0100; 
	if(x==?20'b??1?????001?100?111?) z |= 4'b0100; 
	if(x==?20'b??1??1?0?110??001??1) z |= 4'b1000; 
	if(x==?20'b??11111?0??10?????11) z |= 4'b0100; 
	if(x==?20'b??1?1????101?000?1?1) z |= 4'b1000; 
	if(x==?20'b?1?1111??0?10?????11) z |= 4'b0100; 
	if(x==?20'b??1?1???1?10?000?1?1) z |= 4'b1000; 
	if(x==?20'b?1?????1101?000??1?1) z |= 4'b0100; 
	if(x==?20'b???1?111?11100????1?) z |= 4'b0100; 
	if(x==?20'b????111??0?1?00111??) z |= 4'b1000; 
	if(x==?20'b????1100??01???111??) z |= 4'b1000; 
	if(x==?20'b?1110??????10?1?1?11) z |= 4'b0100; 
	if(x==?20'b?11??10????1001?11??) z |= 4'b0100; 
	if(x==?20'b?111???101??0?0??1?1) z |= 4'b0100; 
	if(x==?20'b?111???1?11100?????1) z |= 4'b0100; 
	if(x==?20'b?1???????100?001111?) z |= 4'b1000; 
	if(x==?20'b?1?????101?1000??1?1) z |= 4'b0100; 
	if(x==?20'b1????11011?0?0??1?1?) z |= 4'b1000; 
	if(x==?20'b?1???1?0?111?000???1) z |= 4'b1000; 
	if(x==?20'b11???110???0??001?1?) z |= 4'b1000; 
	if(x==?20'b111?1?????10?0?0?1?1) z |= 4'b1000; 
	if(x==?20'b1????11011?0??0?1?1?) z |= 4'b1000; 
	if(x==?20'b?11?011?00??0???1?1?) z |= 4'b0100; 
	if(x==?20'b???10111?1??00???11?) z |= 4'b0100; 
	if(x==?20'b?11??110??00???01?1?) z |= 4'b1000; 
	if(x==?20'b?1110??1?1??00???1?1) z |= 4'b0100; 
	if(x==?20'b?1110111?1???1???1??) z |= 4'b0100; 
	if(x==?20'b1???1110??1???00?11?) z |= 4'b1000; 
	if(x==?20'b?1????11111??00???01) z |= 4'b0100; 
	if(x==?20'b111?1??0??1???00?1?1) z |= 4'b1000; 
	if(x==?20'b111?1??0?1???0?0??11) z |= 4'b1000; 
	if(x==?20'b???1011?0?11?0??1?1?) z |= 4'b0100; 
	if(x==?20'b???1011?0?11??0?1?1?) z |= 4'b0100; 
	if(x==?20'b?1??????1100?10?111?) z |= 4'b1000; 
	if(x==?20'b1???11??111??0?0??11) z |= 4'b1000; 
	if(x==?20'b??1?11???111?00???01) z |= 4'b1000; 
	if(x==?20'b?1110??10????00???11) z |= 4'b0100; 
	if(x==?20'b111?1??0???0?00???11) z |= 4'b1000; 
	if(x==?20'b??1?1110??10???0?11?) z |= 4'b1000; 
	if(x==?20'b?1?1???1??110?1?1?11) z |= 4'b0100; 
	if(x==?20'b11??1??0111???0???11) z |= 4'b1000; 
	if(x==?20'b?1110??1??1?0?0???11) z |= 4'b0100; 
	if(x==?20'b111????011????00??11) z |= 4'b1000; 
	if(x==?20'b111?1110??1???1??1??) z |= 4'b1000; 
	if(x==?20'b?11?0???01??000??1?1) z |= 4'b0100; 
	if(x==?20'b??1????10101?00?11??) z |= 4'b0100; 
	if(x==?20'b?11????11011?1???11?) z |= 4'b0100; 
	if(x==?20'b?????111?10?100?11??) z |= 4'b0100; 
	if(x==?20'b??1?1??011???0?11?11) z |= 4'b1000; 
	if(x==?20'b?11?1???1101??1??11?) z |= 4'b1000; 
	if(x==?20'b????11??110??0001?1?) z |= 4'b1000; 
	if(x==?20'b???1??11?1110?0???11) z |= 4'b0100; 
	if(x==?20'b?????1?01110?00?1??1) z |= 4'b1000; 
	if(x==?20'b????1?111?00??0?1?11) z |= 4'b1000; 
	if(x==?20'b?1?10?1?011??0??1??1) z |= 4'b0100; 
	if(x==?20'b?11?11????1111??1??1) z |= 4'b0100; 
	if(x==?20'b?111?111?1??01???1??) z |= 4'b0100; 
	if(x==?20'b??110??1?111?0????11) z |= 4'b0100; 
	if(x==?20'b????0?1?0111?00?1??1) z |= 4'b0100; 
	if(x==?20'b1????11011????001?1?) z |= 4'b1000; 
	if(x==?20'b111?1?????0??000??11) z |= 4'b1000; 
	if(x==?20'b?11????0??10?000?1?1) z |= 4'b1000; 
	if(x==?20'b??1??1??010?000??11?) z |= 4'b0100; 
	if(x==?20'b??110?1?111??00????1) z |= 4'b0100; 
	if(x==?20'b?1110?????1100????11) z |= 4'b0100; 
	if(x==?20'b1?1??1?0?110??0?1??1) z |= 4'b1000; 
	if(x==?20'b????11?100?1?0??1?11) z |= 4'b0100; 
	if(x==?20'b?11?1?11?1??010??1??) z |= 4'b0100; 
	if(x==?20'b?111???10???000???11) z |= 4'b0100; 
	if(x==?20'b111?1??????0?000??11) z |= 4'b1000; 
	if(x==?20'b?111???1?0??000???11) z |= 4'b0100; 
	if(x==?20'b11??1???111???00??11) z |= 4'b1000; 
	if(x==?20'b?11???1111????111??1) z |= 4'b1000; 
	if(x==?20'b??1?????0011?01?111?) z |= 4'b0100; 
	if(x==?20'b??1?0??1011??00?1??1) z |= 4'b0100; 
	if(x==?20'b?1??1??0?110?00?1??1) z |= 4'b1000; 
	if(x==?20'b??1??11011?0???01?1?) z |= 4'b1000; 
	if(x==?20'b?1110?????1?0?1?1?11) z |= 4'b0100; 
	if(x==?20'b??1?11???110?0?11?1?) z |= 4'b1000; 
	if(x==?20'b?1????1??010?000?11?) z |= 4'b1000; 
	if(x==?20'b11???1?0?111?00????1) z |= 4'b1000; 
	if(x==?20'b???1011???1100??1?1?) z |= 4'b0100; 
	if(x==?20'b??????11?011000?1?1?) z |= 4'b0100; 
	if(x==?20'b?????1?0111??000??11) z |= 4'b1000; 
	if(x==?20'b111?1??0?????000??11) z |= 4'b1000; 
	if(x==?20'b?111011?00??????1?1?) z |= 4'b0100; 
	if(x==?20'b111??110??00????1?1?) z |= 4'b1000; 
	if(x==?20'b?11?01?????1010??1?1) z |= 4'b0100; 
	if(x==?20'b?11???101????010?1?1) z |= 4'b1000; 
	if(x==?20'b?1110??1????000???11) z |= 4'b0100; 
	if(x==?20'b?????1??1110?0001??1) z |= 4'b1000; 
	if(x==?20'b?1?1??1?011?00??1??1) z |= 4'b0100; 
	if(x==?20'b??1?0?1?11???00?1?01) z |= 4'b0100; 
	if(x==?20'b??11???1?11100????11) z |= 4'b0100; 
	if(x==?20'b?1??011?0?110???1?1?) z |= 4'b0100; 
	if(x==?20'b????0?1??111000???11) z |= 4'b0100; 
	if(x==?20'b??????1?0111000?1??1) z |= 4'b0100; 
	if(x==?20'b1?????1?11?0??001?11) z |= 4'b1000; 
	if(x==?20'b??11??1?111?000????1) z |= 4'b0100; 
	if(x==?20'b?11?11?1??1??010?1??) z |= 4'b1000; 
	if(x==?20'b111????1???0?0?111?1) z |= 4'b1000; 
	if(x==?20'b1?1??1???110??001??1) z |= 4'b1000; 
	if(x==?20'b1?1?11??11???0?11?1?) z |= 4'b1000; 
	if(x==?20'b1?1?1?10?????000?11?) z |= 4'b1000; 
	if(x==?20'b???1001?010?????11??) z |= 4'b0100; 
	if(x==?20'b????1???11?0?0001?11) z |= 4'b1000; 
	if(x==?20'b??1????1011?000?1??1) z |= 4'b0100; 
	if(x==?20'b?1??1????110?0001??1) z |= 4'b1000; 
	if(x==?20'b?1??101??1??000??11?) z |= 4'b0100; 
	if(x==?20'b?11???1111??11??1?1?) z |= 4'b0100; 
	if(x==?20'b11???1???111?000???1) z |= 4'b1000; 
	if(x==?20'b?1?101?1????000??11?) z |= 4'b0100; 
	if(x==?20'b?1?1??11??111?0?1?1?) z |= 4'b0100; 
	if(x==?20'b?1110???01???00??1?1) z |= 4'b0100; 
	if(x==?20'b?1?1111?0???00????11) z |= 4'b0100; 
	if(x==?20'b?1???0101001????11??) z |= 4'b1100; 
	if(x==?20'b?????1111??0?000??11) z |= 4'b1000; 
	if(x==?20'b1?1??111??0??0?0??11) z |= 4'b1000; 
	if(x==?20'b?1???1?0??11?00?1?01) z |= 4'b1000; 
	if(x==?20'b1???11??110??00?1?1?) z |= 4'b1000; 
	if(x==?20'b??11111?0???0?0???11) z |= 4'b0100; 
	if(x==?20'b?111?11?00??0???1?1?) z |= 4'b0100; 
	if(x==?20'b?1?1111??0??0?0???11) z |= 4'b0100; 
	if(x==?20'b111??11???00???01?1?) z |= 4'b1000; 
	if(x==?20'b????1??011???0001?11) z |= 4'b1000; 
	if(x==?20'b????111?0??1000???11) z |= 4'b0100; 
	if(x==?20'b?11?0?1?111?00?????1) z |= 4'b0100; 
	if(x==?20'b??1???1?11??000?1?01) z |= 4'b0100; 
	if(x==?20'b??1???1?00??111???11) z |= 4'b0100; 
	if(x==?20'b11???111???0?0?0??11) z |= 4'b1000; 
	if(x==?20'b??1??101??1??000?11?) z |= 4'b1000; 
	if(x==?20'b111????0??10?00??1?1) z |= 4'b1000; 
	if(x==?20'b1?1??111???0??00??11) z |= 4'b1000; 
	if(x==?20'b?11??01?1????00111??) z |= 4'b1000; 
	if(x==?20'b1????100?010????11??) z |= 4'b1000; 
	if(x==?20'b???????10?11000?1?11) z |= 4'b0100; 
	if(x==?20'b1?????101????000?111) z |= 4'b1000; 
	if(x==?20'b111????01????0?11?11) z |= 4'b1000; 
	if(x==?20'b??1?11??1100??0?1?1?) z |= 4'b1000; 
	if(x==?20'b??1?11??00??00??1?11) z |= 4'b0100; 
	if(x==?20'b1???11?1??1??000?11?) z |= 4'b1000; 
	if(x==?20'b1?1??11011?0????1?1?) z |= 4'b1000; 
	if(x==?20'b??????11011?000?1?1?) z |= 4'b0100; 
	if(x==?20'b?11??1?0?111??00???1) z |= 4'b1000; 
	if(x==?20'b?1?????1?100???1110?) z |= 4'b1000; 
	if(x==?20'b?1????11??00??001?11) z |= 4'b1000; 
	if(x==?20'b????11???110?0001?1?) z |= 4'b1000; 
	if(x==?20'b????0??1??11000?1?11) z |= 4'b0100; 
	if(x==?20'b???101?????1000??111) z |= 4'b0100; 
	if(x==?20'b?1???1????00?111??11) z |= 4'b1000; 
	if(x==?20'b1????1?0111??00???11) z |= 4'b1000; 
	if(x==?20'b?111????01??000??1?1) z |= 4'b0100; 
	if(x==?20'b11?????011????001?11) z |= 4'b1000; 
	if(x==?20'b???1??11?011?00?1?1?) z |= 4'b0100; 
	if(x==?20'b111?1?1???0??0?0??11) z |= 4'b1000; 
	if(x==?20'b?1???1????11?0001?01) z |= 4'b1000; 
	if(x==?20'b1?1?1???11???0?11?11) z |= 4'b1000; 
	if(x==?20'b?11?1??11????01011??) z |= 4'b1000; 
	if(x==?20'b?11101?????1?10??1?1) z |= 4'b0100; 
	if(x==?20'b111???101????01??1?1) z |= 4'b1000; 
	if(x==?20'b??1?0?1?11?100??1??1) z |= 4'b0100; 
	if(x==?20'b1????1??1110?00?1??1) z |= 4'b1000; 
	if(x==?20'b?11???11111???0???01) z |= 4'b0100; 
	if(x==?20'b?1???1??0?110?1?1?11) z |= 4'b0100; 
	if(x==?20'b?1????110011?0??1?1?) z |= 4'b0100; 
	if(x==?20'b?1?1011?0?11????1?1?) z |= 4'b0100; 
	if(x==?20'b???10?1??111?00???11) z |= 4'b0100; 
	if(x==?20'b?111?1?10???00????11) z |= 4'b0100; 
	if(x==?20'b???1??1?0111?00?1??1) z |= 4'b0100; 
	if(x==?20'b111?1?1????0??00??11) z |= 4'b1000; 
	if(x==?20'b111???????10?000?1?1) z |= 4'b1000; 
	if(x==?20'b?11?11???111?0????01) z |= 4'b1000; 
	if(x==?20'b?11?01??1???010?11??) z |= 4'b0100; 
	if(x==?20'b?111?1?1?0??0?0???11) z |= 4'b0100; 
	if(x==?20'b111?11?1??1??01??1??) z |= 4'b1000; 
	if(x==?20'b????011111??00??1?1?) z |= 4'b0100; 
	if(x==?20'b???????1110??000111?) z |= 4'b1000; 
	if(x==?20'b111???1?1?0???00??11) z |= 4'b1000; 
	if(x==?20'b?1???1?01?11??001??1) z |= 4'b1000; 
	if(x==?20'b?11?11????11??111?1?) z |= 4'b1000; 
	if(x==?20'b?1??0?11111??00????1) z |= 4'b0100; 
	if(x==?20'b????001110????1?11??) z |= 4'b0100; 
	if(x==?20'b1???11??11???0001?1?) z |= 4'b1000; 
	if(x==?20'b11???11?1?00?0??1?1?) z |= 4'b1000; 
	if(x==?20'b11???11?1?00??0?1?1?) z |= 4'b1000; 
	if(x==?20'b111????0?1???000??11) z |= 4'b1000; 
	if(x==?20'b???????111?0?000111?) z |= 4'b1000; 
	if(x==?20'b1?1??11?11?0???01?1?) z |= 4'b1000; 
	if(x==?20'b?11?1???0???010?11?1) z |= 4'b0100; 
	if(x==?20'b??1?11??110???001?1?) z |= 4'b1000; 
	if(x==?20'b??1?11?0?111?00????1) z |= 4'b1000; 
	if(x==?20'b1????1??111??000??11) z |= 4'b1000; 
	if(x==?20'b?1???1?01110?0??1??1) z |= 4'b1000; 
	if(x==?20'b1????1111??0?00???11) z |= 4'b1000; 
	if(x==?20'b?11?????1100??1?111?) z |= 4'b1000; 
	if(x==?20'b?1110?????1?000???11) z |= 4'b0100; 
	if(x==?20'b????1?11??00?00?1?11) z |= 4'b1000; 
	if(x==?20'b??1??1?01110??0?1??1) z |= 4'b1000; 
	if(x==?20'b??1?1???1101?00??1?1) z |= 4'b1000; 
	if(x==?20'b?11?????0011?1??111?) z |= 4'b0100; 
	if(x==?20'b????1110??11??001?1?) z |= 4'b1000; 
	if(x==?20'b?111?1?????1010??1?1) z |= 4'b0100; 
	if(x==?20'b????11?100???00?1?11) z |= 4'b0100; 
	if(x==?20'b?111?1???0?100????11) z |= 4'b0100; 
	if(x==?20'b???1111?0??1?00???11) z |= 4'b0100; 
	if(x==?20'b??11?11?00?1?0??1?1?) z |= 4'b0100; 
	if(x==?20'b111???1?1????010?1?1) z |= 4'b1000; 
	if(x==?20'b????1???0?11000?111?) z |= 4'b0100; 
	if(x==?20'b1?1??11011?????01?1?) z |= 4'b1000; 
	if(x==?20'b?1??0?1?0111?0??1??1) z |= 4'b0100; 
	if(x==?20'b????1????011000?111?) z |= 4'b0100; 
	if(x==?20'b111??1?01????0?0??11) z |= 4'b1000; 
	if(x==?20'b?1?10???1???000?11?1) z |= 4'b0100; 
	if(x==?20'b??11?11?00?1??0?1?1?) z |= 4'b0100; 
	if(x==?20'b??1?0?1?0111??0?1??1) z |= 4'b0100; 
	if(x==?20'b?1?1?11?0?110???1?1?) z |= 4'b0100; 
	if(x==?20'b???1??1??111000???11) z |= 4'b0100; 
	if(x==?20'b?11???10???1?01011??) z |= 4'b1000; 
	if(x==?20'b???1??11??11000?1?1?) z |= 4'b0100; 
	if(x==?20'b11?????01????0001?11) z |= 4'b1000; 
	if(x==?20'b?1110?1????10?0???11) z |= 4'b0100; 
	if(x==?20'b?11??1101?00????1?1?) z |= 4'b1000; 
	if(x==?20'b?1????11111?000????1) z |= 4'b0100; 
	if(x==?20'b1?1????0???1?00011?1) z |= 4'b1000; 
	if(x==?20'b?1?????11011?00??1?1) z |= 4'b0100; 
	if(x==?20'b?11????1???0?01011?1) z |= 4'b1000; 
	if(x==?20'b111????0?1???0?11?11) z |= 4'b1000; 
	if(x==?20'b?1????11?01100??1?1?) z |= 4'b0100; 
	if(x==?20'b?11?0?????110?1?1?11) z |= 4'b0100; 
	if(x==?20'b?1???1?0111??0?0??11) z |= 4'b1000; 
	if(x==?20'b???1??11011??00?1?1?) z |= 4'b0100; 
	if(x==?20'b?1?1011???110???1?1?) z |= 4'b0100; 
	if(x==?20'b????11??00?1?00?1?11) z |= 4'b0100; 
	if(x==?20'b??1??1?0111???00??11) z |= 4'b1000; 
	if(x==?20'b??110??????1000?1?11) z |= 4'b0100; 
	if(x==?20'b???10??1??11?00?1?11) z |= 4'b0100; 
	if(x==?20'b??1?11???111?000???1) z |= 4'b1000; 
	if(x==?20'b?1???1??1110?0?01??1) z |= 4'b1000; 
	if(x==?20'b?11?011?00?1????1?1?) z |= 4'b0100; 
	if(x==?20'b??1??1??1110??001??1) z |= 4'b1000; 
	if(x==?20'b1???1???11???0001?11) z |= 4'b1000; 
	if(x==?20'b?1??0?1??11100????11) z |= 4'b0100; 
	if(x==?20'b?1????1?011100??1??1) z |= 4'b0100; 
	if(x==?20'b??1???10??00?00??111) z |= 4'b1000; 
	if(x==?20'b??1?0?1??1110?0???11) z |= 4'b0100; 
	if(x==?20'b??1???1?01110?0?1??1) z |= 4'b0100; 
	if(x==?20'b?1??01??00???00??111) z |= 4'b0100; 
	if(x==?20'b111??1??111??0?0???1) z |= 4'b1000; 
	if(x==?20'b?11???1111???11?1??1) z |= 4'b1000; 
	if(x==?20'b1???1?0??100??0?11??) z |= 4'b1000; 
	if(x==?20'b11???11?1??0??001?1?) z |= 4'b1000; 
	if(x==?20'b???1011111???0??1?1?) z |= 4'b0100; 
	if(x==?20'b??1??1111?0??0?0??11) z |= 4'b1000; 
	if(x==?20'b????111?111??000??1?) z |= 4'b1000; 
	if(x==?20'b?11??11?1?00???01?1?) z |= 4'b1000; 
	if(x==?20'b?11?0011?1???0??1?1?) z |= 4'b0100; 
	if(x==?20'b???1?0?1001??0??11??) z |= 4'b0100; 
	if(x==?20'b?11?0011?1????0?1?1?) z |= 4'b0100; 
	if(x==?20'b?111??1??1110?0????1) z |= 4'b0100; 
	if(x==?20'b?1111???0????10?11?1) z |= 4'b0100; 
	if(x==?20'b?1???1111??0?0?0??11) z |= 4'b1000; 
	if(x==?20'b??1??1111??0??00??11) z |= 4'b1000; 
	if(x==?20'b?11?1100??1???0?1?1?) z |= 4'b1000; 
	if(x==?20'b111?1???11???0?0??11) z |= 4'b1000; 
	if(x==?20'b1?1?11??110???0?1?1?) z |= 4'b1000; 
	if(x==?20'b???1???1??11000?1?11) z |= 4'b0100; 
	if(x==?20'b?1??111?0??100????11) z |= 4'b0100; 
	if(x==?20'b?11?11????11?11?1??1) z |= 4'b0100; 
	if(x==?20'b??1?1??011????001?11) z |= 4'b1000; 
	if(x==?20'b??1?111?0??10?0???11) z |= 4'b0100; 
	if(x==?20'b?11??11?00?10???1?1?) z |= 4'b0100; 
	if(x==?20'b?1??111??0?10?0???11) z |= 4'b0100; 
	if(x==?20'b1???1110??11??0?1?1?) z |= 4'b1000; 
	if(x==?20'b?????111?111000???1?) z |= 4'b0100; 
	if(x==?20'b111?1???1??0?00???11) z |= 4'b1000; 
	if(x==?20'b??1???1???00?000?111) z |= 4'b1000; 
	if(x==?20'b???111???11?000?1?1?) z |= 4'b0100; 
	if(x==?20'b?1???1??00??000??111) z |= 4'b0100; 
	if(x==?20'b1?????11?11??0001?1?) z |= 4'b1000; 
	if(x==?20'b???1?11111??00??1?1?) z |= 4'b0100; 
	if(x==?20'b111?1??01????00???11) z |= 4'b1000; 
	if(x==?20'b????0111?1??000??11?) z |= 4'b0100; 
	if(x==?20'b?111???10??1?00???11) z |= 4'b0100; 
	if(x==?20'b?1?1??11111??00????1) z |= 4'b0100; 
	if(x==?20'b??1?0?1?11??000?1??1) z |= 4'b0100; 
	if(x==?20'b????1110??1??000?11?) z |= 4'b1000; 
	if(x==?20'b??1???1?11?0?0?11?11) z |= 4'b1000; 
	if(x==?20'b??1?11???110??001?1?) z |= 4'b1000; 
	if(x==?20'b?1?1??11?011?0??1?1?) z |= 4'b0100; 
	if(x==?20'b?111???1??110?0???11) z |= 4'b0100; 
	if(x==?20'b11?????0?1???0001?11) z |= 4'b1000; 
	if(x==?20'b1?1??1?0111???0???11) z |= 4'b1000; 
	if(x==?20'b?1?1??11?011??0?1?1?) z |= 4'b0100; 
	if(x==?20'b1?1??10?110????0?1??) z |= 4'b1000; 
	if(x==?20'b1?1?11???111?00????1) z |= 4'b1000; 
	if(x==?20'b1?1??1??1110??0?1??1) z |= 4'b1000; 
	if(x==?20'b??110?????1?000?1?11) z |= 4'b0100; 
	if(x==?20'b1???111???11??001?1?) z |= 4'b1000; 
	if(x==?20'b?1110??1???1?00???11) z |= 4'b0100; 
	if(x==?20'b?1??1??0111??00???11) z |= 4'b1000; 
	if(x==?20'b?1?10?1??111?0????11) z |= 4'b0100; 
	if(x==?20'b?1?1??1?0111?0??1??1) z |= 4'b0100; 
	if(x==?20'b???10??1101??1???11?) z |= 4'b0100; 
	if(x==?20'b?11?01101??1?0??1?1?) z |= 4'b1100; 
	if(x==?20'b1???110?10?????011??) z |= 4'b1000; 
	if(x==?20'b?11?01101??1??0?1?1?) z |= 4'b1100; 
	if(x==?20'b?11??????100?10?111?) z |= 4'b1000; 
	if(x==?20'b?1??1???1110?00?1??1) z |= 4'b1000; 
	if(x==?20'b?11???1?111??00???01) z |= 4'b0100; 
	if(x==?20'b111???1???0??000??11) z |= 4'b1000; 
	if(x==?20'b?1???1?0??11?0001??1) z |= 4'b1000; 
	if(x==?20'b?11??110110??0??1???) z |= 4'b1000; 
	if(x==?20'b?11??110110???0?1???) z |= 4'b1000; 
	if(x==?20'b??1?1???001??1??110?) z |= 4'b0100; 
	if(x==?20'b?11?0?11111???0????1) z |= 4'b0100; 
	if(x==?20'b1?1??1111?0??0????11) z |= 4'b1000; 
	if(x==?20'b1???111?111??00???1?) z |= 4'b1000; 
	if(x==?20'b111?1???1????000??11) z |= 4'b1000; 
	if(x==?20'b1?1?11??11????001?1?) z |= 4'b1000; 
	if(x==?20'b?1?1?01??0110????1??) z |= 4'b0100; 
	if(x==?20'b111??11?1?00????1?1?) z |= 4'b1000; 
	if(x==?20'b?111?1???0??000???11) z |= 4'b0100; 
	if(x==?20'b?11???1111???11?1?1?) z |= 4'b0100; 
	if(x==?20'b111?1???111??00????1) z |= 4'b1000; 
	if(x==?20'b?1??0?1?011??00?1??1) z |= 4'b0100; 
	if(x==?20'b1???1??0?101??1??11?) z |= 4'b1000; 
	if(x==?20'b?????11011???0001?1?) z |= 4'b1000; 
	if(x==?20'b??1?0??1?111?00???11) z |= 4'b0100; 
	if(x==?20'b??1????10111?00?1??1) z |= 4'b0100; 
	if(x==?20'b??1???1??101?000?11?) z |= 4'b1000; 
	if(x==?20'b?11?11?0?111?0?????1) z |= 4'b1000; 
	if(x==?20'b?1????1??101?000?11?) z |= 4'b1000; 
	if(x==?20'b11???1??111??0?0??11) z |= 4'b1000; 
	if(x==?20'b?111??????110?1?1?11) z |= 4'b0100; 
	if(x==?20'b?11??1???111?00???01) z |= 4'b1000; 
	if(x==?20'b??1??1??101?000??11?) z |= 4'b0100; 
	if(x==?20'b?1???1??101?000??11?) z |= 4'b0100; 
	if(x==?20'b11???1111??0?0????11) z |= 4'b1000; 
	if(x==?20'b1?1??1??111???00??11) z |= 4'b1000; 
	if(x==?20'b?11????011???0001??1) z |= 4'b1000; 
	if(x==?20'b1?1??1111??0??0???11) z |= 4'b1000; 
	if(x==?20'b??1???1?1?10?000?11?) z |= 4'b1000; 
	if(x==?20'b?1????1?1?10?000?11?) z |= 4'b1000; 
	if(x==?20'b??1??1?0?110?00?1??1) z |= 4'b1000; 
	if(x==?20'b??1?1?11??00??0?1?11) z |= 4'b1000; 
	if(x==?20'b?1??1?11??00??0?1?11) z |= 4'b1000; 
	if(x==?20'b??1?11?100???0??1?11) z |= 4'b0100; 
	if(x==?20'b?1??11?100???0??1?11) z |= 4'b0100; 
	if(x==?20'b?1?1111?0??1?0????11) z |= 4'b0100; 
	if(x==?20'b??1??1??01?1000??11?) z |= 4'b0100; 
	if(x==?20'b?1???1??01?1000??11?) z |= 4'b0100; 
	if(x==?20'b??1?11?100????0?1?11) z |= 4'b0100; 
	if(x==?20'b??11111?0??1??0???11) z |= 4'b0100; 
	if(x==?20'b??11011??1??00??1?1?) z |= 4'b0100; 
	if(x==?20'b?111?11?00?1????1?1?) z |= 4'b0100; 
	if(x==?20'b?1?1111??0?1??0???11) z |= 4'b0100; 
	if(x==?20'b?1?????1?100??1?110?) z |= 4'b1000; 
	if(x==?20'b?1110???1???0?0?11?1) z |= 4'b0100; 
	if(x==?20'b??1?1???001???1?110?) z |= 4'b0100; 
	if(x==?20'b?111???1???1000???11) z |= 4'b0100; 
	if(x==?20'b???1?111?111?00???1?) z |= 4'b0100; 
	if(x==?20'b?1??1???111??000??11) z |= 4'b1000; 
	if(x==?20'b1???1???1100???011??) z |= 4'b1000; 
	if(x==?20'b?1?1??1??11100????11) z |= 4'b0100; 
	if(x==?20'b?11?11????11?11?1?1?) z |= 4'b1000; 
	if(x==?20'b?????11?1011?1??01??) z |= 4'b0100; 
	if(x==?20'b11????1?1??1?0?11?11) z |= 4'b1000; 
	if(x==?20'b??11??1??1110?0???11) z |= 4'b0100; 
	if(x==?20'b1????111?1???0001??1) z |= 4'b1000; 
	if(x==?20'b1?1?1?1?1????000?11?) z |= 4'b1000; 
	if(x==?20'b?11?011??011?0??1???) z |= 4'b0100; 
	if(x==?20'b?111???1?111?00????1) z |= 4'b0100; 
	if(x==?20'b?11???????00?0001?11) z |= 4'b1000; 
	if(x==?20'b?11????011???0?11?11) z |= 4'b1000; 
	if(x==?20'b11???110???0?00?1?1?) z |= 4'b1000; 
	if(x==?20'b?11?011??011??0?1???) z |= 4'b0100; 
	if(x==?20'b?????11?1101??1?01??) z |= 4'b1000; 
	if(x==?20'b??1???111?00??0?1?11) z |= 4'b1000; 
	if(x==?20'b????011???11000?1?1?) z |= 4'b0100; 
	if(x==?20'b?1????111?00??0?1?11) z |= 4'b1000; 
	if(x==?20'b?11??1???0?10?1?1?11) z |= 4'b0100; 
	if(x==?20'b111????01?????001?11) z |= 4'b1000; 
	if(x==?20'b111?1???11????0011??) z |= 4'b1000; 
	if(x==?20'b1????01?1100????11??) z |= 4'b1000; 
	if(x==?20'b111????0???1?0?011?1) z |= 4'b1000; 
	if(x==?20'b???10011?10?????11??) z |= 4'b0100; 
	if(x==?20'b?11?0?????11000?1??1) z |= 4'b0100; 
	if(x==?20'b?11???11111?0?0????1) z |= 4'b0100; 
	if(x==?20'b???10111?1???00??11?) z |= 4'b0100; 
	if(x==?20'b1???1110??1??00??11?) z |= 4'b1000; 
	if(x==?20'b??1?11??00?1?0??1?11) z |= 4'b0100; 
	if(x==?20'b?1????1?011?000?1??1) z |= 4'b0100; 
	if(x==?20'b?1??11??00?1?0??1?11) z |= 4'b0100; 
	if(x==?20'b?1110??1?1???00??1?1) z |= 4'b0100; 
	if(x==?20'b??1????1?111000???11) z |= 4'b0100; 
	if(x==?20'b111?1??0??1??00??1?1) z |= 4'b1000; 
	if(x==?20'b111?111?1????0?0??1?) z |= 4'b1000; 
	if(x==?20'b???1?11?1?1?000?1??1) z |= 4'b0100; 
	if(x==?20'b??????1?11?0?0001?11) z |= 4'b1000; 
	if(x==?20'b?1?1011?????000??11?) z |= 4'b0100; 
	if(x==?20'b?11?11???111?0?0???1) z |= 4'b1000; 
	if(x==?20'b1???1100?01?????11??) z |= 4'b1000; 
	if(x==?20'b111?1?1?1??0??0???11) z |= 4'b1000; 
	if(x==?20'b?1?1?1?1???1000??11?) z |= 4'b0100; 
	if(x==?20'b??1??1???110?0001??1) z |= 4'b1000; 
	if(x==?20'b???1???100110???11??) z |= 4'b0100; 
	if(x==?20'b1?1?1???11????001?11) z |= 4'b1000; 
	if(x==?20'b1?1?111?1????0?0??11) z |= 4'b1000; 
	if(x==?20'b1?1???101????0?0111?) z |= 4'b1000; 
	if(x==?20'b??1???11?0??111???11) z |= 4'b0100; 
	if(x==?20'b?111???1??1100??11??) z |= 4'b0100; 
	if(x==?20'b???1?10?0011????11??) z |= 4'b0100; 
	if(x==?20'b11???1111?????00??11) z |= 4'b1000; 
	if(x==?20'b?1??1?11??0???001?11) z |= 4'b1000; 
	if(x==?20'b111????011???00???11) z |= 4'b1000; 
	if(x==?20'b?111?1?10??1?0????11) z |= 4'b0100; 
	if(x==?20'b?1??11????0??111??11) z |= 4'b1000; 
	if(x==?20'b?11?01101?1??0??1?1?) z |= 4'b1100; 
	if(x==?20'b?????1??0?11000?1?11) z |= 4'b0100; 
	if(x==?20'b?1??111?111??0?0??1?) z |= 4'b1000; 
	if(x==?20'b?111?111???10?0???1?) z |= 4'b0100; 
	if(x==?20'b?11?01101?1???0?1?1?) z |= 4'b1100; 
	if(x==?20'b??1?111?111???00??1?) z |= 4'b1000; 
	if(x==?20'b?1??111?0???000???11) z |= 4'b0100; 
	if(x==?20'b??1?11?1?0??00??1?11) z |= 4'b0100; 
	if(x==?20'b??11111????100????11) z |= 4'b0100; 
	if(x==?20'b?11?0110?1?1?0??1?1?) z |= 4'b1100; 
	if(x==?20'b???1?111?1??000??11?) z |= 4'b0100; 
	if(x==?20'b?1?101?????10?0?111?) z |= 4'b0100; 
	if(x==?20'b?11?0110?1?1??0?1?1?) z |= 4'b1100; 
	if(x==?20'b??11011?????000?1?1?) z |= 4'b0100; 
	if(x==?20'b11????1?11???0001??1) z |= 4'b1000; 
	if(x==?20'b11???110?????0001?1?) z |= 4'b1000; 
	if(x==?20'b?1?1?111???10?0???11) z |= 4'b0100; 
	if(x==?20'b?111???1?1??000??1?1) z |= 4'b0100; 
	if(x==?20'b1????11011???00?1?1?) z |= 4'b1000; 
	if(x==?20'b?111?111?1???10??1??) z |= 4'b0100; 
	if(x==?20'b?11??1111??0???0??11) z |= 4'b1000; 
	if(x==?20'b??1??111???0?000??11) z |= 4'b1000; 
	if(x==?20'b111?1?????1??000?1?1) z |= 4'b1000; 
	if(x==?20'b?11?111?0??10?????11) z |= 4'b0100; 
	if(x==?20'b?1???111?11100????1?) z |= 4'b0100; 
	if(x==?20'b?1110?????11?00???11) z |= 4'b0100; 
	if(x==?20'b?1??????11?0?0001?11) z |= 4'b1000; 
	if(x==?20'b??1??111?1110?0???1?) z |= 4'b0100; 
	if(x==?20'b?11??1?1???1010?11??) z |= 4'b0100; 
	if(x==?20'b11??1???111??00???11) z |= 4'b1000; 
	if(x==?20'b??1??11011?0?0??1?1?) z |= 4'b1000; 
	if(x==?20'b?11??110???0??001?1?) z |= 4'b1000; 
	if(x==?20'b??1??0111100????11??) z |= 4'b1100; 
	if(x==?20'b??1??11011?0??0?1?1?) z |= 4'b1000; 
	if(x==?20'b???1?01?0?01?0??11??) z |= 4'b0100; 
	if(x==?20'b111?????11???000??11) z |= 4'b1000; 
	if(x==?20'b1????10?10?0??0?11??) z |= 4'b1000; 
	if(x==?20'b?1?????011???0001?11) z |= 4'b1000; 
	if(x==?20'b?1??0111?1??00???11?) z |= 4'b0100; 
	if(x==?20'b???1011???11?00?1?1?) z |= 4'b0100; 
	if(x==?20'b??11?1????11000?1??1) z |= 4'b0100; 
	if(x==?20'b????0?1110??0?1?11??) z |= 4'b0100; 
	if(x==?20'b111??11?110??0??1???) z |= 4'b1000; 
	if(x==?20'b????110?1?01??1?11??) z |= 4'b1000; 
	if(x==?20'b111??11?110???0?1???) z |= 4'b1000; 
	if(x==?20'b??1?????0?11000?1?11) z |= 4'b0100; 
	if(x==?20'b??1?1110??1???00?11?) z |= 4'b1000; 
	if(x==?20'b????11?0??01??1011??) z |= 4'b1000; 
	if(x==?20'b??11?1???0??000?1?11) z |= 4'b0100; 
	if(x==?20'b?1?1??1?011??00?1??1) z |= 4'b0100; 
	if(x==?20'b?1??011?0?11?0??1?1?) z |= 4'b0100; 
	if(x==?20'b111????0?1????001?11) z |= 4'b1000; 
	if(x==?20'b1????11?11???0001?1?) z |= 4'b1000; 
	if(x==?20'b???1?11?11??000?1?1?) z |= 4'b0100; 
	if(x==?20'b??11???1?111?00???11) z |= 4'b0100; 
	if(x==?20'b1?1??10??10??0?0?1??) z |= 4'b1000; 
	if(x==?20'b?1??011?0?11??0?1?1?) z |= 4'b0100; 
	if(x==?20'b?1??110?0011????11??) z |= 4'b1100; 
	if(x==?20'b??1?11??111??0?0??11) z |= 4'b1000; 
	if(x==?20'b1?1??1???110?00?1??1) z |= 4'b1000; 
	if(x==?20'b?111??????11000???11) z |= 4'b0100; 
	if(x==?20'b??1?0?????11000?1?11) z |= 4'b0100; 
	if(x==?20'b?11?1??0111???0???11) z |= 4'b1000; 
	if(x==?20'b??1?0??1010??1???11?) z |= 4'b0100; 
	if(x==?20'b?1?1?01??01?0?0??1??) z |= 4'b0100; 
	if(x==?20'b????0??10??101???111) z |= 4'b0100; 
	if(x==?20'b?111?111?1??00????1?) z |= 4'b0100; 
	if(x==?20'b?????100?1???10011??) z |= 4'b1000; 
	if(x==?20'b?111?11??011?0??1???) z |= 4'b0100; 
	if(x==?20'b111?????11???0?11?11) z |= 4'b1000; 
	if(x==?20'b?111?11??011??0?1???) z |= 4'b0100; 
	if(x==?20'b????1??01??0??10?111) z |= 4'b1000; 
	if(x==?20'b111?111???1???00??1?) z |= 4'b1000; 
	if(x==?20'b???1?1??0?11?00?1?11) z |= 4'b0100; 
	if(x==?20'b1????11???11?0001?1?) z |= 4'b1000; 
	if(x==?20'b???1?11???11000?1?1?) z |= 4'b0100; 
	if(x==?20'b1?1?111?111???0???1?) z |= 4'b1000; 
	if(x==?20'b?1????11?1110?0???11) z |= 4'b0100; 
	if(x==?20'b?1?1111?0????00???11) z |= 4'b0100; 
	if(x==?20'b?111?1??1???0?1?1?11) z |= 4'b0100; 
	if(x==?20'b?111?11?00???0??1?1?) z |= 4'b0100; 
	if(x==?20'b111??11???00?0??1?1?) z |= 4'b1000; 
	if(x==?20'b?111?11?00????0?1?1?) z |= 4'b0100; 
	if(x==?20'b111??11???00??0?1?1?) z |= 4'b1000; 
	if(x==?20'b?11?0??1?111?0????11) z |= 4'b0100; 
	if(x==?20'b??1??11011????001?1?) z |= 4'b1000; 
	if(x==?20'b?11?0?1?111??00????1) z |= 4'b0100; 
	if(x==?20'b1?1??111???0?00???11) z |= 4'b1000; 
	if(x==?20'b????001???1?001?11??) z |= 4'b0100; 
	if(x==?20'b?1?1?111?111?0????1?) z |= 4'b0100; 
	if(x==?20'b?11?1???111???00??11) z |= 4'b1000; 
	if(x==?20'b?1??1??0?010??1??11?) z |= 4'b1000; 
	if(x==?20'b?11??1?0?111?00????1) z |= 4'b1000; 
	if(x==?20'b?1??011???1100??1?1?) z |= 4'b0100; 
	if(x==?20'b???1?01????1010?11??) z |= 4'b0100; 
	if(x==?20'b??1??11011?1?00?1?1?) z |= 4'b1100; 
	if(x==?20'b111????0?????0001?11) z |= 4'b1000; 
	if(x==?20'b11??1?10?1?0???0?1??) z |= 4'b1000; 
	if(x==?20'b?1110?1?11???0??1??1) z |= 4'b0100; 
	if(x==?20'b?1??011?1?11?00?1?1?) z |= 4'b1100; 
	if(x==?20'b1????10?1????01011??) z |= 4'b1000; 
	if(x==?20'b?11????1?11100????11) z |= 4'b0100; 
	if(x==?20'b??1?0?1?11?1?00?1??1) z |= 4'b0100; 
	if(x==?20'b??1101?10?1?0????1??) z |= 4'b0100; 
	if(x==?20'b?1????1???00?101?1?1) z |= 4'b1000; 
	if(x==?20'b??1???1?11?0??001?11) z |= 4'b1000; 
	if(x==?20'b111?111??????000??1?) z |= 4'b1000; 
	if(x==?20'b?11???1?111?000????1) z |= 4'b0100; 
	if(x==?20'b111?1?1????0?00???11) z |= 4'b1000; 
	if(x==?20'b??1??1??00??101??1?1) z |= 4'b0100; 
	if(x==?20'b?111?1?10????00???11) z |= 4'b0100; 
	if(x==?20'b?111?111????000???1?) z |= 4'b0100; 
	if(x==?20'b111???1?1?0??00???11) z |= 4'b1000; 
	if(x==?20'b?1???1?01?11?00?1??1) z |= 4'b1000; 
	if(x==?20'b????011111???00?1?1?) z |= 4'b0100; 
	if(x==?20'b??11111?????000???11) z |= 4'b0100; 
	if(x==?20'b??110?????11?00?1?11) z |= 4'b0100; 
	if(x==?20'b??1??01?0101?0???1??) z |= 4'b0100; 
	if(x==?20'b11???111?????000??11) z |= 4'b1000; 
	if(x==?20'b1?1??11?11?0?0??1?1?) z |= 4'b1000; 
	if(x==?20'b?11??1???111?000???1) z |= 4'b1000; 
	if(x==?20'b111??11????0??001?1?) z |= 4'b1000; 
	if(x==?20'b?????011?011??1?11??) z |= 4'b0100; 
	if(x==?20'b1?1??11?11?0??0?1?1?) z |= 4'b1000; 
	if(x==?20'b111??1?0??11??0?1??1) z |= 4'b1000; 
	if(x==?20'b?1??1?11?11???001?1?) z |= 4'b1000; 
	if(x==?20'b1?1?1?1?1?1??1?1?1??) z |= 4'b1000; 
	if(x==?20'b??1?11?1?11?00??1?1?) z |= 4'b0100; 
	if(x==?20'b?11?111?0???0?0???11) z |= 4'b0100; 
	if(x==?20'b11??????11???0001?11) z |= 4'b1000; 
	if(x==?20'b?1???10?1010??0??1??) z |= 4'b1000; 
	if(x==?20'b????1110??11?00?1?1?) z |= 4'b1000; 
	if(x==?20'b1?1?1?1??1?1?1?1?1??) z |= 4'b1000; 
	if(x==?20'b?111??1?11??00??1??1) z |= 4'b0100; 
	if(x==?20'b1?1??1?11?1??1?1?1??) z |= 4'b1000; 
	if(x==?20'b1?1??11011???0??1?1?) z |= 4'b1000; 
	if(x==?20'b1????10??1?0?0?0?11?) z |= 4'b1000; 
	if(x==?20'b???1?01?0?1?0?0??11?) z |= 4'b0100; 
	if(x==?20'b?111?1???0?1?00???11) z |= 4'b0100; 
	if(x==?20'b?1?11?1??1?11?1??1??) z |= 4'b0100; 
	if(x==?20'b?11??111???0?0?0??11) z |= 4'b1000; 
	if(x==?20'b1?1??11011????0?1?1?) z |= 4'b1000; 
	if(x==?20'b??1???1?11?1000?1??1) z |= 4'b0100; 
	if(x==?20'b?1?1?1?11?1?1?1??1??) z |= 4'b0100; 
	if(x==?20'b?1?1?11?0?11?0??1?1?) z |= 4'b0100; 
	if(x==?20'b??1???101????000?111) z |= 4'b1000; 
	if(x==?20'b?1?1?11?0?11??0?1?1?) z |= 4'b0100; 
	if(x==?20'b?11?1???001??0??111?) z |= 4'b0100; 
	if(x==?20'b?1?1?1?1?1?11?1??1??) z |= 4'b0100; 
	if(x==?20'b?1???1??1?11?0001??1) z |= 4'b1000; 
	if(x==?20'b?????11111??000?1?1?) z |= 4'b0100; 
	if(x==?20'b??11??????11000?1?11) z |= 4'b0100; 
	if(x==?20'b??1?11?1??1??000?11?) z |= 4'b1000; 
	if(x==?20'b???1???10??101???111) z |= 4'b0100; 
	if(x==?20'b11????1?1??1??001?11) z |= 4'b1000; 
	if(x==?20'b?1?1011???11?0??1?1?) z |= 4'b0100; 
	if(x==?20'b??1??1?0111??00???11) z |= 4'b1000; 
	if(x==?20'b?11????011????001?11) z |= 4'b1000; 
	if(x==?20'b?1??01?????1000??111) z |= 4'b0100; 
	if(x==?20'b?1?1011???11??0?1?1?) z |= 4'b0100; 
	if(x==?20'b111??1????11??001??1) z |= 4'b1000; 
	if(x==?20'b1???1???1??0??10?111) z |= 4'b1000; 
	if(x==?20'b?1??1?0?1?00??0?11??) z |= 4'b1000; 
	if(x==?20'b?????1?0??01?10011??) z |= 4'b1000; 
	if(x==?20'b??1??1??1110?00?1??1) z |= 4'b1000; 
	if(x==?20'b????111???11?0001?1?) z |= 4'b1000; 
	if(x==?20'b?1??1?101010?????1??) z |= 4'b1000; 
	if(x==?20'b?1??0?1??111?00???11) z |= 4'b0100; 
	if(x==?20'b1?1??11?11????001?1?) z |= 4'b1000; 
	if(x==?20'b?1????1?0111?00?1??1) z |= 4'b0100; 
	if(x==?20'b??1?01?10101?????1??) z |= 4'b0100; 
	if(x==?20'b1???1?0???0???00111?) z |= 4'b1000; 
	if(x==?20'b??1??0?1?001?0??11??) z |= 4'b0100; 
	if(x==?20'b????11?0??01?0?111??) z |= 4'b1000; 
	if(x==?20'b?1??1?111?0???0?1?11) z |= 4'b1000; 
	if(x==?20'b11???11?1??0?00?1?1?) z |= 4'b1000; 
	if(x==?20'b???1?0?1?0??00??111?) z |= 4'b0100; 
	if(x==?20'b??1?11??11???0001?1?) z |= 4'b1000; 
	if(x==?20'b??11?11??1?100??1?1?) z |= 4'b0100; 
	if(x==?20'b?11??11?1?00?0??1?1?) z |= 4'b1000; 
	if(x==?20'b?11??11?1?00??0?1?1?) z |= 4'b1000; 
	if(x==?20'b1???11?0???0??001??1) z |= 4'b1000; 
	if(x==?20'b?1?1?11???1100??1?1?) z |= 4'b0100; 
	if(x==?20'b??1??1??111??000??11) z |= 4'b1000; 
	if(x==?20'b????1???1??0?101?111) z |= 4'b1000; 
	if(x==?20'b??1?11?1?0?1?0??1?11) z |= 4'b0100; 
	if(x==?20'b?11??11?00?1?0??1?1?) z |= 4'b0100; 
	if(x==?20'b?11??11?00?1??0?1?1?) z |= 4'b0100; 
	if(x==?20'b1?1?1?1??11??1?1?1??) z |= 4'b1000; 
	if(x==?20'b?1????1??111000???11) z |= 4'b0100; 
	if(x==?20'b?1?11?1??11?1?1??1??) z |= 4'b0100; 
	if(x==?20'b???????10??1101??111) z |= 4'b0100; 
	if(x==?20'b?1????11??11000?1?1?) z |= 4'b0100; 
	if(x==?20'b?11????01????0001?11) z |= 4'b1000; 
	if(x==?20'b1?1??1?1?11??1?1?1??) z |= 4'b1000; 
	if(x==?20'b11??1????100???011??) z |= 4'b1000; 
	if(x==?20'b?1?1?1?1?11?1?1??1??) z |= 4'b0100; 
	if(x==?20'b???1?11111???00?1?1?) z |= 4'b0100; 
	if(x==?20'b???10?1?0?01?0??11??) z |= 4'b0100; 
	if(x==?20'b1????1?010?0??0?11??) z |= 4'b1000; 
	if(x==?20'b?1????11011??00?1?1?) z |= 4'b0100; 
	if(x==?20'b????11?01?01??1?11??) z |= 4'b1000; 
	if(x==?20'b??1?0110010?????11??) z |= 4'b1100; 
	if(x==?20'b11???11?1????0001?1?) z |= 4'b1000; 
	if(x==?20'b?11?0??????1000?1?11) z |= 4'b0100; 
	if(x==?20'b?1??0??1??11?00?1?11) z |= 4'b0100; 
	if(x==?20'b1?1??10?110??0???1??) z |= 4'b1000; 
	if(x==?20'b??11???1001?0???11??) z |= 4'b0100; 
	if(x==?20'b????1100?1???10?11??) z |= 4'b1000; 
	if(x==?20'b??1?1???11???0001?11) z |= 4'b1000; 
	if(x==?20'b1???111???11?00?1?1?) z |= 4'b1000; 
	if(x==?20'b????001???1?100?11??) z |= 4'b0110; 
	if(x==?20'b???1111?00??0?????11) z |= 4'b0100; 
	if(x==?20'b?1??1?1011????10?1??) z |= 4'b1000; 
	if(x==?20'b??11?1???0?1?00?1?11) z |= 4'b0100; 
	if(x==?20'b??11?11????1000?1?1?) z |= 4'b0100; 
	if(x==?20'b?1???1111????000??11) z |= 4'b1000; 
	if(x==?20'b??1?1?0??100??0?11??) z |= 4'b1000; 
	if(x==?20'b1?1??10??010????11??) z |= 4'b1000; 
	if(x==?20'b?11??11?1??0??001?1?) z |= 4'b1000; 
	if(x==?20'b????11???010??0111??) z |= 4'b1000; 
	if(x==?20'b1????111??00???0??11) z |= 4'b1000; 
	if(x==?20'b?1??0110?010????11??) z |= 4'b1100; 
	if(x==?20'b??1?011111???0??1?1?) z |= 4'b0100; 
	if(x==?20'b?1??011111???0??1?1?) z |= 4'b0100; 
	if(x==?20'b??1?01?1??1101???1??) z |= 4'b0100; 
	if(x==?20'b?????100?1???00111??) z |= 4'b1001; 
	if(x==?20'b??1?111????1000???11) z |= 4'b0100; 
	if(x==?20'b?1???0?1001??0??11??) z |= 4'b0100; 
	if(x==?20'b?1?1?01??011??0??1??) z |= 4'b0100; 
	if(x==?20'b???1?011??01??0?11??) z |= 4'b0100; 
	if(x==?20'b????0011??1??01?11??) z |= 4'b0100; 
	if(x==?20'b????11??1?01??1011??) z |= 4'b1000; 
	if(x==?20'b1?1??1??111??00???11) z |= 4'b1000; 
	if(x==?20'b111?????11????001?11) z |= 4'b1000; 
	if(x==?20'b?1?????1??11000?1?11) z |= 4'b0100; 
	if(x==?20'b????110??1???10011??) z |= 4'b1000; 
	if(x==?20'b??1?1110??11??0?1?1?) z |= 4'b1000; 
	if(x==?20'b?1??1110??11??0?1?1?) z |= 4'b1000; 
	if(x==?20'b1???111?1??0??00???1) z |= 4'b1000; 
	if(x==?20'b??11011??1???00?1?1?) z |= 4'b0100; 
	if(x==?20'b1???1???1100?0??11??) z |= 4'b1000; 
	if(x==?20'b?1??11???11??0001?1?) z |= 4'b1000; 
	if(x==?20'b??1?11???11?000?1?1?) z |= 4'b0100; 
	if(x==?20'b?1??11???11?000?1?1?) z |= 4'b0100; 
	if(x==?20'b11??1?1?1010?????1??) z |= 4'b1000; 
	if(x==?20'b??1???11?11??0001?1?) z |= 4'b1000; 
	if(x==?20'b?1????11?11??0001?1?) z |= 4'b1000; 
	if(x==?20'b?1?1??1??111?00???11) z |= 4'b0100; 
	if(x==?20'b??1???11?11?000?1?1?) z |= 4'b0100; 
	if(x==?20'b??11?1?10101?????1??) z |= 4'b0100; 
	if(x==?20'b??1??11111??00??1?1?) z |= 4'b0100; 
	if(x==?20'b?1???11111??00??1?1?) z |= 4'b0100; 
	if(x==?20'b111?1???11???00?11??) z |= 4'b1000; 
	if(x==?20'b???1?1110??100?????1) z |= 4'b0100; 
	if(x==?20'b??1?0??1?1??101??11?) z |= 4'b0100; 
	if(x==?20'b?1??1??0??1??101?11?) z |= 4'b1000; 
	if(x==?20'b11????1????1?0001?11) z |= 4'b1000; 
	if(x==?20'b?11????0?1???0001?11) z |= 4'b1000; 
	if(x==?20'b?????011??1?001?11??) z |= 4'b0100; 
	if(x==?20'b?1110??????1?00?1?11) z |= 4'b0100; 
	if(x==?20'b?11?0?????1?000?1?11) z |= 4'b0100; 
	if(x==?20'b??1?111???11??001?1?) z |= 4'b1000; 
	if(x==?20'b?1??111???11??001?1?) z |= 4'b1000; 
	if(x==?20'b???1???10011??0?11??) z |= 4'b0100; 
	if(x==?20'b??11?11??1??000?1?1?) z |= 4'b0100; 
	if(x==?20'b??1?0??1101??1???11?) z |= 4'b0100; 
	if(x==?20'b?1??0??1101??1???11?) z |= 4'b0100; 
	if(x==?20'b??1??11?11?100??1?1?) z |= 4'b0100; 
	if(x==?20'b??1?110?10?????011??) z |= 4'b1000; 
	if(x==?20'b??1??1??00??010??1?1) z |= 4'b0100; 
	if(x==?20'b11???1111????00???11) z |= 4'b1000; 
	if(x==?20'b?111???1??11?00?11??) z |= 4'b0100; 
	if(x==?20'b?1??1?11??0??00?1?11) z |= 4'b1000; 
	if(x==?20'b????11?01??0??001??1) z |= 4'b1000; 
	if(x==?20'b11???11???1??0001?1?) z |= 4'b1000; 
	if(x==?20'b?1?1?01?0???0?0??11?) z |= 4'b0100; 
	if(x==?20'b?1???11?1?11??001?1?) z |= 4'b1000; 
	if(x==?20'b????0?11?011??1?11??) z |= 4'b0100; 
	if(x==?20'b??1?11?1?0???00?1?11) z |= 4'b0100; 
	if(x==?20'b??11111????1?00???11) z |= 4'b0100; 
	if(x==?20'b1?1??10????0?0?0?11?) z |= 4'b1000; 
	if(x==?20'b??1?1??0?101??1??11?) z |= 4'b1000; 
	if(x==?20'b?1??1??0?101??1??11?) z |= 4'b1000; 
	if(x==?20'b?11??1??111??0?0??11) z |= 4'b1000; 
	if(x==?20'b?1????1???00?010?1?1) z |= 4'b1000; 
	if(x==?20'b1?1?11??1?10???0?1??) z |= 4'b1000; 
	if(x==?20'b?111???????1000?1?11) z |= 4'b0100; 
	if(x==?20'b?1?1???1??11?00?1?11) z |= 4'b0100; 
	if(x==?20'b????0?1110???10?11??) z |= 4'b0100; 
	if(x==?20'b??1???1?00??11??1?11) z |= 4'b0100; 
	if(x==?20'b?1?1??1101?10????1??) z |= 4'b0100; 
	if(x==?20'b?11?011??1??00??1?1?) z |= 4'b0100; 
	if(x==?20'b???1011????10?1?1??1) z |= 4'b0100; 
	if(x==?20'b??1?1???1100???011??) z |= 4'b1000; 
	if(x==?20'b1?1??110?1?0???0?1??) z |= 4'b1000; 
	if(x==?20'b?1??1???1100???011??) z |= 4'b1000; 
	if(x==?20'b???1?0?1????100?111?) z |= 4'b0100; 
	if(x==?20'b?111??1?11?1?0??1??1) z |= 4'b0100; 
	if(x==?20'b?1?1011?0?1?0????1??) z |= 4'b0100; 
	if(x==?20'b?11???1?1??1?0?11?11) z |= 4'b1000; 
	if(x==?20'b11??11??110????01???) z |= 4'b1000; 
	if(x==?20'b?11???1??1110?0???11) z |= 4'b0100; 
	if(x==?20'b11??1?1?11????10?1??) z |= 4'b1000; 
	if(x==?20'b?1??110?101???0??1??) z |= 4'b1000; 
	if(x==?20'b?1??0011?10?????11??) z |= 4'b0100; 
	if(x==?20'b111??1??1?11??0?1??1) z |= 4'b1000; 
	if(x==?20'b??1??011?101?0???1??) z |= 4'b0100; 
	if(x==?20'b??11?1?1??1101???1??) z |= 4'b0100; 
	if(x==?20'b1???1?0??????001111?) z |= 4'b1000; 
	if(x==?20'b?1??0111?1???00??11?) z |= 4'b0100; 
	if(x==?20'b1????1101?0????011??) z |= 4'b1000; 
	if(x==?20'b?1??1??0100???0?11??) z |= 4'b1000; 
	if(x==?20'b?????1?01?01?10?11??) z |= 4'b1000; 
	if(x==?20'b??1?1110??1??00??11?) z |= 4'b1000; 
	if(x==?20'b??????11?0110?1?11??) z |= 4'b0100; 
	if(x==?20'b??1?1100?01?????11??) z |= 4'b1000; 
	if(x==?20'b11??1??011?0????1??1) z |= 4'b1000; 
	if(x==?20'b??1????100110???11??) z |= 4'b0100; 
	if(x==?20'b?1?????100110???11??) z |= 4'b0100; 
	if(x==?20'b??????1110??010?11??) z |= 4'b0100; 
	if(x==?20'b?????1111?00???0??11) z |= 4'b1000; 
	if(x==?20'b11??1?10???0???0?11?) z |= 4'b1000; 
	if(x==?20'b??1101?10???0????11?) z |= 4'b0100; 
	if(x==?20'b??1?01?1??1?010??1??) z |= 4'b0100; 
	if(x==?20'b?1110?????1??00?1?11) z |= 4'b0100; 
	if(x==?20'b??11??11?0110???1???) z |= 4'b0100; 
	if(x==?20'b1?1??11?1?1??1?1?1??) z |= 4'b1000; 
	if(x==?20'b???1011??0?10???11??) z |= 4'b0100; 
	if(x==?20'b?11?1??11?1??00?1?11) z |= 4'b1100; 
	if(x==?20'b?1??1?10?1???010?1??) z |= 4'b1000; 
	if(x==?20'b????111?00?10?????11) z |= 4'b0100; 
	if(x==?20'b?1???1????00??111?11) z |= 4'b1000; 
	if(x==?20'b?11??1111?????00??11) z |= 4'b1000; 
	if(x==?20'b11??11????00???01?1?) z |= 4'b1000; 
	if(x==?20'b????0??10??1?10??111) z |= 4'b0100; 
	if(x==?20'b??11??1100??0???1?1?) z |= 4'b0100; 
	if(x==?20'b?11?1??1?1?1?00?1?11) z |= 4'b1100; 
	if(x==?20'b?1?1?11??1?11?1??1??) z |= 4'b0100; 
	if(x==?20'b?111?111?1???00???1?) z |= 4'b0100; 
	if(x==?20'b?????10??10??000?11?) z |= 4'b1000; 
	if(x==?20'b????1??01??0?01??111) z |= 4'b1000; 
	if(x==?20'b111?111???1??00???1?) z |= 4'b1000; 
	if(x==?20'b?11?111????100????11) z |= 4'b0100; 
	if(x==?20'b??110??10?11????1??1) z |= 4'b0100; 
	if(x==?20'b?1???111?1??000??11?) z |= 4'b0100; 
	if(x==?20'b?11???1?11???0001??1) z |= 4'b1000; 
	if(x==?20'b?11?011?????000?1?1?) z |= 4'b0100; 
	if(x==?20'b?11??110?????0001?1?) z |= 4'b1000; 
	if(x==?20'b?????01??01?000??11?) z |= 4'b0100; 
	if(x==?20'b????11????01?01011??) z |= 4'b1000; 
	if(x==?20'b1???111???0??000???1) z |= 4'b1000; 
	if(x==?20'b111??????1???0001?11) z |= 4'b1000; 
	if(x==?20'b?11??010???1?10?11??) z |= 4'b1100; 
	if(x==?20'b??1?0??101??00???1?1) z |= 4'b0100; 
	if(x==?20'b11??1???11?0???01??1) z |= 4'b1000; 
	if(x==?20'b???1?1110???000????1) z |= 4'b0100; 
	if(x==?20'b1???111????0?000???1) z |= 4'b1000; 
	if(x==?20'b???1?111?0??000????1) z |= 4'b0100; 
	if(x==?20'b?11?010?1????01?11??) z |= 4'b1100; 
	if(x==?20'b?111??????1?000?1?11) z |= 4'b0100; 
	if(x==?20'b?11?01100??0?????11?) z |= 4'b1100; 
	if(x==?20'b?11?1???111??00???11) z |= 4'b1000; 
	if(x==?20'b??????11010??01?11??) z |= 4'b0100; 
	if(x==?20'b1?1?1?10?10???0??1??) z |= 4'b1000; 
	if(x==?20'b???1011???1?0?1?1??1) z |= 4'b0100; 
	if(x==?20'b?1??1??0??10??00?1?1) z |= 4'b1000; 
	if(x==?20'b11??1??011?????01??1) z |= 4'b1000; 
	if(x==?20'b?1???01?0?01?0??11??) z |= 4'b0100; 
	if(x==?20'b???????10??1010??111) z |= 4'b0100; 
	if(x==?20'b??1??10?10?0??0?11??) z |= 4'b1000; 
	if(x==?20'b1???1?1011?????0?11?) z |= 4'b1000; 
	if(x==?20'b?11??1????11000?1??1) z |= 4'b0100; 
	if(x==?20'b11??1?10?1?0?0???1??) z |= 4'b1000; 
	if(x==?20'b????1???1??0?010?111) z |= 4'b1000; 
	if(x==?20'b?????011??1?100?11??) z |= 4'b0100; 
	if(x==?20'b??11???10?110???1??1) z |= 4'b0100; 
	if(x==?20'b????11?0??10?10?11??) z |= 4'b1000; 
	if(x==?20'b111???1????1??001?11) z |= 4'b1000; 
	if(x==?20'b?11??1???0??000?1?11) z |= 4'b0100; 
	if(x==?20'b??1??11?11???0001?1?) z |= 4'b1000; 
	if(x==?20'b??1??11?11??000?1?1?) z |= 4'b0100; 
	if(x==?20'b?1???11?11??000?1?1?) z |= 4'b0100; 
	if(x==?20'b?1?101?1?01??0???1??) z |= 4'b0100; 
	if(x==?20'b?11????1?111?00???11) z |= 4'b0100; 
	if(x==?20'b????110??1???00111??) z |= 4'b1000; 
	if(x==?20'b??1101?10?1???0??1??) z |= 4'b0100; 
	if(x==?20'b??11??11011?0???1???) z |= 4'b0100; 
	if(x==?20'b?111?11??1??00??1?1?) z |= 4'b0100; 
	if(x==?20'b11??11???110???01???) z |= 4'b1000; 
	if(x==?20'b?1?????0?100?1??111?) z |= 4'b1000; 
	if(x==?20'b??????1?01010?0??11?) z |= 4'b0100; 
	if(x==?20'b??110??1??110???1??1) z |= 4'b0100; 
	if(x==?20'b1?1??1?0?010????11??) z |= 4'b1000; 
	if(x==?20'b?????1??1010?0?0?11?) z |= 4'b1000; 
	if(x==?20'b??1?0???001??1??111?) z |= 4'b0100; 
	if(x==?20'b????11?0???0?0001??1) z |= 4'b1000; 
	if(x==?20'b???101?1??110????11?) z |= 4'b0100; 
	if(x==?20'b111??11????0?00?1?1?) z |= 4'b1000; 
	if(x==?20'b?1??1?11?11??00?1?1?) z |= 4'b1000; 
	if(x==?20'b?1???1??0?11?00?1?11) z |= 4'b0100; 
	if(x==?20'b??1??11???11?0001?1?) z |= 4'b1000; 
	if(x==?20'b?1???11???11?0001?1?) z |= 4'b1000; 
	if(x==?20'b?1???11???11000?1?1?) z |= 4'b0100; 
	if(x==?20'b??1?11?1?11??00?1?1?) z |= 4'b0100; 
	if(x==?20'b??1??10?1?0??0?011??) z |= 4'b1000; 
	if(x==?20'b?1?1?11??11?1?1??1??) z |= 4'b0100; 
	if(x==?20'b?1?1?011?10?????11??) z |= 4'b0100; 
	if(x==?20'b????11????10?10011??) z |= 4'b1000; 
	if(x==?20'b?111??1?11???00?1??1) z |= 4'b0100; 
	if(x==?20'b?1?????0?100??1?111?) z |= 4'b1000; 
	if(x==?20'b??11?11??11?11??1???) z |= 4'b0100; 
	if(x==?20'b????0?1??011?01?11??) z |= 4'b0100; 
	if(x==?20'b1?1?110??01?????11??) z |= 4'b1000; 
	if(x==?20'b1????1101????0?11??1) z |= 4'b1000; 
	if(x==?20'b??110??101???0???1?1) z |= 4'b0100; 
	if(x==?20'b??1?0???001???1?111?) z |= 4'b0100; 
	if(x==?20'b?11?0??11?00????1?11) z |= 4'b1100; 
	if(x==?20'b?1??1????100?0?011??) z |= 4'b1000; 
	if(x==?20'b??????110?1?001?11??) z |= 4'b0100; 
	if(x==?20'b??11?1?1??1?010??1??) z |= 4'b0100; 
	if(x==?20'b?????0?1???1100?111?) z |= 4'b0100; 
	if(x==?20'b11??1?1??1???010?1??) z |= 4'b1000; 
	if(x==?20'b??110??1????0?1?1?11) z |= 4'b0100; 
	if(x==?20'b11??1??0??10??0??1?1) z |= 4'b1000; 
	if(x==?20'b??1??01????1010?11??) z |= 4'b0100; 
	if(x==?20'b?1???01????1010?11??) z |= 4'b0100; 
	if(x==?20'b???1???10??1?10??111) z |= 4'b0100; 
	if(x==?20'b?11?1?10?1?0???0?1??) z |= 4'b1000; 
	if(x==?20'b111??1????11?00?1??1) z |= 4'b1000; 
	if(x==?20'b111???1???0??00?1?11) z |= 4'b1000; 
	if(x==?20'b??1?0??1?1??010??11?) z |= 4'b0100; 
	if(x==?20'b???10?11011?????1?1?) z |= 4'b0100; 
	if(x==?20'b1???1???1??0?01??111) z |= 4'b1000; 
	if(x==?20'b??1????1001?0?0?11??) z |= 4'b0100; 
	if(x==?20'b??1??11111?1?0??1?1?) z |= 4'b0100; 
	if(x==?20'b?1???10?1????01011??) z |= 4'b1000; 
	if(x==?20'b?1??1?101??0???0?11?) z |= 4'b1000; 
	if(x==?20'b1???11?0?110????1?1?) z |= 4'b1000; 
	if(x==?20'b?1??111?1?11??0?1?1?) z |= 4'b1000; 
	if(x==?20'b?11?01?10?1?0????1??) z |= 4'b0100; 
	if(x==?20'b?111?1???0???00?1?11) z |= 4'b0100; 
	if(x==?20'b111??11??????0001?1?) z |= 4'b1000; 
	if(x==?20'b?111?11?????000?1?1?) z |= 4'b0100; 
	if(x==?20'b1?1??11?11???00?1?1?) z |= 4'b1000; 
	if(x==?20'b????111?00??0?0???11) z |= 4'b0100; 
	if(x==?20'b?????111??00?0?0??11) z |= 4'b1000; 
	if(x==?20'b11???11??11???111???) z |= 4'b1000; 
	if(x==?20'b??11???101??00???1?1) z |= 4'b0100; 
	if(x==?20'b????1?0?1????001111?) z |= 4'b1010; 
	if(x==?20'b?11?111?????000???11) z |= 4'b0100; 
	if(x==?20'b1?1??10?1?0???0??11?) z |= 4'b1000; 
	if(x==?20'b??1?01?10??10????11?) z |= 4'b0100; 
	if(x==?20'b?11?0?????11?00?1?11) z |= 4'b0100; 
	if(x==?20'b???10?11?1??00??1??1) z |= 4'b0100; 
	if(x==?20'b?1??1??0??1??010?11?) z |= 4'b1000; 
	if(x==?20'b?11??111?????000??11) z |= 4'b1000; 
	if(x==?20'b??11?11??1?1?00?1?1?) z |= 4'b0100; 
	if(x==?20'b11??1?????10??00?1?1) z |= 4'b1000; 
	if(x==?20'b1???11?0???0?00?1??1) z |= 4'b1000; 
	if(x==?20'b????111?1?0??000???1) z |= 4'b1000; 
	if(x==?20'b?11?????11???0001?11) z |= 4'b1000; 
	if(x==?20'b?1?1?01??0?1?0???11?) z |= 4'b0100; 
	if(x==?20'b?1?1?11???11?00?1?1?) z |= 4'b0100; 
	if(x==?20'b?11?1?100??0?0???11?) z |= 4'b1100; 
	if(x==?20'b??1??10??1?0?0?0?11?) z |= 4'b1000; 
	if(x==?20'b????111?1??0?000???1) z |= 4'b1000; 
	if(x==?20'b?1???01?0?1?0?0??11?) z |= 4'b0100; 
	if(x==?20'b?11?01?10??0??0??11?) z |= 4'b1100; 
	if(x==?20'b??1???1?00???11?1?11) z |= 4'b0100; 
	if(x==?20'b1?1??110?101?????1??) z |= 4'b1000; 
	if(x==?20'b111?1??01??0??????11) z |= 4'b1000; 
	if(x==?20'b?1???1????00?11?1?11) z |= 4'b1000; 
	if(x==?20'b?1?1?1110???00?????1) z |= 4'b0100; 
	if(x==?20'b1?1??1101?10?????1??) z |= 4'b1000; 
	if(x==?20'b?1?1011?01?1?????1??) z |= 4'b0100; 
	if(x==?20'b1?1?111????0??00???1) z |= 4'b1000; 
	if(x==?20'b?????1110??1000????1) z |= 4'b0100; 
	if(x==?20'b11??1????100?0??11??) z |= 4'b1000; 
	if(x==?20'b?????111?0?1000????1) z |= 4'b0100; 
	if(x==?20'b?11???????11000?1?11) z |= 4'b0100; 
	if(x==?20'b1????110?1???0?11??1) z |= 4'b1000; 
	if(x==?20'b?1?????10??101???111) z |= 4'b0100; 
	if(x==?20'b?11???1?1??1??001?11) z |= 4'b1000; 
	if(x==?20'b????011???110?1?1??1) z |= 4'b0100; 
	if(x==?20'b?1110??10??1??????11) z |= 4'b0100; 
	if(x==?20'b1???1?10?1???0?0?11?) z |= 4'b1000; 
	if(x==?20'b??1??1100110????11??) z |= 4'b1100; 
	if(x==?20'b??11??1?011?0?0??1??) z |= 4'b0100; 
	if(x==?20'b??1?1???1??0??10?111) z |= 4'b1000; 
	if(x==?20'b??1101??1???10??11??) z |= 4'b0100; 
	if(x==?20'b?111??1?0101?????1??) z |= 4'b0100; 
	if(x==?20'b??11???1001???0?11??) z |= 4'b0100; 
	if(x==?20'b11??1?101??0?????11?) z |= 4'b1000; 
	if(x==?20'b11???1???110?0?0?1??) z |= 4'b1000; 
	if(x==?20'b1?1??10?1????0?0?11?) z |= 4'b1000; 
	if(x==?20'b111??1??1010?????1??) z |= 4'b1000; 
	if(x==?20'b?1??1?1011???01??1??) z |= 4'b1000; 
	if(x==?20'b???1111?00????0???11) z |= 4'b0100; 
	if(x==?20'b11??11??1?00????1?1?) z |= 4'b1000; 
	if(x==?20'b???101?1??1?0?0??11?) z |= 4'b0100; 
	if(x==?20'b1?1??110?????1?01??1) z |= 4'b1000; 
	if(x==?20'b1????111??00?0????11) z |= 4'b1000; 
	if(x==?20'b?1???10???0??000?11?) z |= 4'b1000; 
	if(x==?20'b?11101?1??1??1???1??) z |= 4'b0100; 
	if(x==?20'b??1??01??0??000??11?) z |= 4'b0100; 
	if(x==?20'b?1?1?01????10?0??11?) z |= 4'b0100; 
	if(x==?20'b??1101?10??1?????11?) z |= 4'b0100; 
	if(x==?20'b?11??11??1?100??1?1?) z |= 4'b0100; 
	if(x==?20'b??1?01?1??11?10??1??) z |= 4'b0100; 
	if(x==?20'b?111???1?1???00?1?11) z |= 4'b0100; 
	if(x==?20'b??1?1?0??????100111?) z |= 4'b1000; 
	if(x==?20'b?????1?0?10??000?11?) z |= 4'b1000; 
	if(x==?20'b??1?11?0???0??001??1) z |= 4'b1000; 
	if(x==?20'b????11??1?01?01?11??) z |= 4'b1000; 
	if(x==?20'b??11??1100?1????1?1?) z |= 4'b0100; 
	if(x==?20'b1???111?11???0?0???1) z |= 4'b1000; 
	if(x==?20'b11????10???1??0111??) z |= 4'b1000; 
	if(x==?20'b????0?1??01?000??11?) z |= 4'b0100; 
	if(x==?20'b11??11?01??0????1?1?) z |= 4'b1000; 
	if(x==?20'b1?1?1????10???0011??) z |= 4'b1000; 
	if(x==?20'b?1?1011?????0?1?1??1) z |= 4'b0100; 
	if(x==?20'b??????1101??100?11??) z |= 4'b0100; 
	if(x==?20'b11??1?1?1??0???0?11?) z |= 4'b1000; 
	if(x==?20'b1???111?1??0?00????1) z |= 4'b1000; 
	if(x==?20'b?1??1?1?11???010?1??) z |= 4'b1000; 
	if(x==?20'b1?1?11??1110?????1??) z |= 4'b1000; 
	if(x==?20'b11??1????1?0??0011??) z |= 4'b1000; 
	if(x==?20'b11?????1???0??0111?1) z |= 4'b1000; 
	if(x==?20'b?1???0?1????001?111?) z |= 4'b0100; 
	if(x==?20'b11??1?101??????0?11?) z |= 4'b1000; 
	if(x==?20'b??11???10?1?00??11??) z |= 4'b0100; 
	if(x==?20'b?1?1011?0???0????11?) z |= 4'b0100; 
	if(x==?20'b?11?1????100???011??) z |= 4'b1000; 
	if(x==?20'b?1?1???1?01?00??11??) z |= 4'b0100; 
	if(x==?20'b??1??11111???00?1?1?) z |= 4'b0100; 
	if(x==?20'b???1?1110??1?00????1) z |= 4'b0100; 
	if(x==?20'b??11?1?10??10????11?) z |= 4'b0100; 
	if(x==?20'b??1??1?1??11010??1??) z |= 4'b0100; 
	if(x==?20'b?111??????11?00?1?11) z |= 4'b0100; 
	if(x==?20'b?1?1??110111?????1??) z |= 4'b0100; 
	if(x==?20'b1?1??110???0???0?11?) z |= 4'b1000; 
	if(x==?20'b???1?111??110?0????1) z |= 4'b0100; 
	if(x==?20'b11??1??0?????0?11?11) z |= 4'b1000; 
	if(x==?20'b?11??11?1????0001?1?) z |= 4'b1000; 
	if(x==?20'b?????11???01?10011??) z |= 4'b1000; 
	if(x==?20'b???1111??0??00????11) z |= 4'b0100; 
	if(x==?20'b1????111??0???00??11) z |= 4'b1000; 
	if(x==?20'b?11????1001?0???11??) z |= 4'b0100; 
	if(x==?20'b1???111????0?0?0??11) z |= 4'b1000; 
	if(x==?20'b????11????10?00111??) z |= 4'b1000; 
	if(x==?20'b?1??1?10???0?0?0?11?) z |= 4'b1000; 
	if(x==?20'b???1?1110???0?0???11) z |= 4'b0100; 
	if(x==?20'b11??1?101??????011??) z |= 4'b1000; 
	if(x==?20'b?1??111???11?00?1?1?) z |= 4'b1000; 
	if(x==?20'b?????11?10??001?11??) z |= 4'b0100; 
	if(x==?20'b??1?01?10???0?0??11?) z |= 4'b0100; 
	if(x==?20'b??1101?1???10????11?) z |= 4'b0100; 
	if(x==?20'b11??11??1110????1???) z |= 4'b1000; 
	if(x==?20'b?1??111?00??0?????11) z |= 4'b0100; 
	if(x==?20'b?11??1???0?1?00?1?11) z |= 4'b0100; 
	if(x==?20'b?11??11????1000?1?1?) z |= 4'b0100; 
	if(x==?20'b1???11?0111???????11) z |= 4'b1000; 
	if(x==?20'b1?1?1?1?110???0??1??) z |= 4'b1000; 
	if(x==?20'b??1??111??00???0??11) z |= 4'b1000; 
	if(x==?20'b????11?01??0?00?1??1) z |= 4'b1000; 
	if(x==?20'b??11011?011?????1???) z |= 4'b0100; 
	if(x==?20'b??11??110111????1???) z |= 4'b0100; 
	if(x==?20'b1???111?1????000???1) z |= 4'b1000; 
	if(x==?20'b11????1?11?0???01??1) z |= 4'b1000; 
	if(x==?20'b????1?1101??00???11?) z |= 4'b0100; 
	if(x==?20'b????0?11?1?100??1??1) z |= 4'b0100; 
	if(x==?20'b??1101?1???10???11??) z |= 4'b0100; 
	if(x==?20'b11???110?110????1???) z |= 4'b1000; 
	if(x==?20'b????11??1?10?10?11??) z |= 4'b1000; 
	if(x==?20'b?1???011??01??0?11??) z |= 4'b0100; 
	if(x==?20'b???10?11?111??????11) z |= 4'b0100; 
	if(x==?20'b???1?11???110?1?1??1) z |= 4'b0100; 
	if(x==?20'b??1?1111010?????11??) z |= 4'b1100; 
	if(x==?20'b??????101??0??00?111) z |= 4'b1000; 
	if(x==?20'b1?1?11??1?10?0???1??) z |= 4'b1000; 
	if(x==?20'b??1???11111??0????01) z |= 4'b0100; 
	if(x==?20'b??????111?00?00?1?11) z |= 4'b1100; 
	if(x==?20'b?1?101?101??????11??) z |= 4'b0100; 
	if(x==?20'b????01??0??100???111) z |= 4'b0100; 
	if(x==?20'b?1?1??1101?1??0??1??) z |= 4'b0100; 
	if(x==?20'b??1?111?1??0??00???1) z |= 4'b1000; 
	if(x==?20'b??????11?011?10?11??) z |= 4'b0100; 
	if(x==?20'b11???11??11??11?1???) z |= 4'b1000; 
	if(x==?20'b??11?1??0?110???1??1) z |= 4'b0100; 
	if(x==?20'b???1?111???1000????1) z |= 4'b0100; 
	if(x==?20'b????11?1??10??00?11?) z |= 4'b1000; 
	if(x==?20'b??11?11??11??11?1???) z |= 4'b0100; 
	if(x==?20'b??1?1???1100?0??11??) z |= 4'b1000; 
	if(x==?20'b1?1??110?1?0?0???1??) z |= 4'b1000; 
	if(x==?20'b?1??1???1100?0??11??) z |= 4'b1000; 
	if(x==?20'b?1????101????10011??) z |= 4'b1000; 
	if(x==?20'b?11?1?1?1010?????1??) z |= 4'b1000; 
	if(x==?20'b1?1?1?10??10????11??) z |= 4'b1000; 
	if(x==?20'b11??11??110??0??1???) z |= 4'b1000; 
	if(x==?20'b11??11??110???0?1???) z |= 4'b1000; 
	if(x==?20'b11??1?1?11???01??1??) z |= 4'b1000; 
	if(x==?20'b?1?1011?0?1???0??1??) z |= 4'b0100; 
	if(x==?20'b?????11011???0?11??1) z |= 4'b1000; 
	if(x==?20'b?1??11???111??0???01) z |= 4'b1000; 
	if(x==?20'b1?1????0?1???000?1?1) z |= 4'b1000; 
	if(x==?20'b?11??1?10101?????1??) z |= 4'b0100; 
	if(x==?20'b?1?1?1?1?011?0???1??) z |= 4'b0100; 
	if(x==?20'b????0?1???110?1?1?11) z |= 4'b0100; 
	if(x==?20'b1????1101?????001??1) z |= 4'b1000; 
	if(x==?20'b?1???1110??100?????1) z |= 4'b0100; 
	if(x==?20'b111?1????100????11??) z |= 4'b1000; 
	if(x==?20'b?1?10?????1?000??1?1) z |= 4'b0100; 
	if(x==?20'b??????110?11?01?11??) z |= 4'b0100; 
	if(x==?20'b??11?1?1??11?10??1??) z |= 4'b0100; 
	if(x==?20'b?11???1????1?0001?11) z |= 4'b1000; 
	if(x==?20'b1?1?1?10?1?????0?11?) z |= 4'b1000; 
	if(x==?20'b?1???1111010????11??) z |= 4'b1100; 
	if(x==?20'b?111???1001?????11??) z |= 4'b0100; 
	if(x==?20'b111?111???00??????1?) z |= 4'b1000; 
	if(x==?20'b??1??1101????1?01??1) z |= 4'b1000; 
	if(x==?20'b?????1111?00?0????11) z |= 4'b1000; 
	if(x==?20'b?1?????1???0?10011?1) z |= 4'b1000; 
	if(x==?20'b11??1?10???0?0???11?) z |= 4'b1000; 
	if(x==?20'b??1????10011??0?11??) z |= 4'b0100; 
	if(x==?20'b1?1?1?10???0??0??11?) z |= 4'b1000; 
	if(x==?20'b?1?????10011??0?11??) z |= 4'b0100; 
	if(x==?20'b?1?101?10????0???11?) z |= 4'b0100; 
	if(x==?20'b11??11???10????01?1?) z |= 4'b1000; 
	if(x==?20'b?111?11100????????1?) z |= 4'b0100; 
	if(x==?20'b??1101?10?????0??11?) z |= 4'b0100; 
	if(x==?20'b??11??11?011?0??1???) z |= 4'b0100; 
	if(x==?20'b?11??11??1??000?1?1?) z |= 4'b0100; 
	if(x==?20'b??11??11?011??0?1???) z |= 4'b0100; 
	if(x==?20'b??1?111001?1????11??) z |= 4'b1100; 
	if(x==?20'b??1?1???0???001?11?1) z |= 4'b0100; 
	if(x==?20'b??1?01?????1001?11??) z |= 4'b0100; 
	if(x==?20'b?1?101?1??1?0????11?) z |= 4'b0100; 
	if(x==?20'b?11??1111????00???11) z |= 4'b1000; 
	if(x==?20'b11??11????00?0??1?1?) z |= 4'b1000; 
	if(x==?20'b????111?00?1??0???11) z |= 4'b0100; 
	if(x==?20'b11??11????00??0?1?1?) z |= 4'b1000; 
	if(x==?20'b11??1??11????10?11??) z |= 4'b1000; 
	if(x==?20'b??11??1100???0??1?1?) z |= 4'b0100; 
	if(x==?20'b?11??11???1??0001?1?) z |= 4'b1000; 
	if(x==?20'b??11??1100????0?1?1?) z |= 4'b0100; 
	if(x==?20'b???1011????1?10?11??) z |= 4'b0100; 
	if(x==?20'b1???1?101??????0111?) z |= 4'b1000; 
	if(x==?20'b??11??11?01?0???1?1?) z |= 4'b0100; 
	if(x==?20'b?11?111????1?00???11) z |= 4'b0100; 
	if(x==?20'b1????1101????01?11??) z |= 4'b1000; 
	if(x==?20'b???11?1101???0???11?) z |= 4'b0100; 
	if(x==?20'b??11???1???10?1?1?11) z |= 4'b0100; 
	if(x==?20'b11??1???11?0?0??1??1) z |= 4'b1000; 
	if(x==?20'b11??1???11?0??0?1??1) z |= 4'b1000; 
	if(x==?20'b??1?0??101???00??1?1) z |= 4'b0100; 
	if(x==?20'b11??1?1????0?0?0?11?) z |= 4'b1000; 
	if(x==?20'b?1??011????10?1?1??1) z |= 4'b0100; 
	if(x==?20'b?11?11??110????01???) z |= 4'b1000; 
	if(x==?20'b1???11?1??10??0??11?) z |= 4'b1000; 
	if(x==?20'b??11?1?10???0?0??11?) z |= 4'b0100; 
	if(x==?20'b???101?1???10???111?) z |= 4'b0100; 
	if(x==?20'b?11?1?1?11????10?1??) z |= 4'b1000; 
	if(x==?20'b1?1????011?0????1?11) z |= 4'b1000; 
	if(x==?20'b?1??1??0??10?00??1?1) z |= 4'b1000; 
	if(x==?20'b11??1??011???0??1??1) z |= 4'b1000; 
	if(x==?20'b11??1??011????0?1??1) z |= 4'b1000; 
	if(x==?20'b??111??1???1?01?11??) z |= 4'b0100; 
	if(x==?20'b1???1?1011???0???11?) z |= 4'b1000; 
	if(x==?20'b?????1111?0???00??11) z |= 4'b1000; 
	if(x==?20'b?11??1?1??1101???1??) z |= 4'b0100; 
	if(x==?20'b????111?1??0?0?0??11) z |= 4'b1000; 
	if(x==?20'b11????10???1?10?11??) z |= 4'b1000; 
	if(x==?20'b??11???10?11?0??1??1) z |= 4'b0100; 
	if(x==?20'b??11???10?11??0?1??1) z |= 4'b0100; 
	if(x==?20'b??11111??0??0?????11) z |= 4'b0100; 
	if(x==?20'b1????110?1????001??1) z |= 4'b1000; 
	if(x==?20'b11???111??0????0??11) z |= 4'b1000; 
	if(x==?20'b?1?10???0?11????1?11) z |= 4'b0100; 
	if(x==?20'b?????11?10??100?11??) z |= 4'b0100; 
	if(x==?20'b??1??1101??0???011??) z |= 4'b1000; 
	if(x==?20'b????111??0?100????11) z |= 4'b0100; 
	if(x==?20'b??1101??1????01?11??) z |= 4'b0100; 
	if(x==?20'b?11?1??011?0????1??1) z |= 4'b1000; 
	if(x==?20'b1?????1?1??0??00?111) z |= 4'b1000; 
	if(x==?20'b?11?1?10???0???0?11?) z |= 4'b1000; 
	if(x==?20'b?11?01?10???0????11?) z |= 4'b0100; 
	if(x==?20'b??11??11011??0??1???) z |= 4'b0100; 
	if(x==?20'b?????1110??10?0???11) z |= 4'b0100; 
	if(x==?20'b??1????101??000??1?1) z |= 4'b0100; 
	if(x==?20'b?11???11?0110???1???) z |= 4'b0100; 
	if(x==?20'b??11??11011???0?1???) z |= 4'b0100; 
	if(x==?20'b11??11???110?0??1???) z |= 4'b1000; 
	if(x==?20'b?1??011??0?10???11??) z |= 4'b0100; 
	if(x==?20'b1???111???1??0?11??1) z |= 4'b1000; 
	if(x==?20'b1?1?1???1?????10111?) z |= 4'b1000; 
	if(x==?20'b???1?1??0??100???111) z |= 4'b0100; 
	if(x==?20'b??110??1??11?0??1??1) z |= 4'b0100; 
	if(x==?20'b11??11???110??0?1???) z |= 4'b1000; 
	if(x==?20'b?111?11??1???00?1?1?) z |= 4'b0100; 
	if(x==?20'b????0?11?1??000?1??1) z |= 4'b0100; 
	if(x==?20'b??110??1??11??0?1??1) z |= 4'b0100; 
	if(x==?20'b?11?11????00???01?1?) z |= 4'b1000; 
	if(x==?20'b?1???1?0??0??000?11?) z |= 4'b1000; 
	if(x==?20'b??111???0????01?11?1) z |= 4'b0100; 
	if(x==?20'b??1?0?1??0??000??11?) z |= 4'b0100; 
	if(x==?20'b?11???1100??0???1?1?) z |= 4'b0100; 
	if(x==?20'b?1??1?????10?000?1?1) z |= 4'b1000; 
	if(x==?20'b??1??110?1???1?01??1) z |= 4'b1000; 
	if(x==?20'b1????11?11???0?11??1) z |= 4'b1000; 
	if(x==?20'b11??1???11????001??1) z |= 4'b1000; 
	if(x==?20'b11??111?1????0?0???1) z |= 4'b1000; 
	if(x==?20'b???101?1??11??0??11?) z |= 4'b0100; 
	if(x==?20'b1???1?1?11???0?0?11?) z |= 4'b1000; 
	if(x==?20'b???1??1???110?1?1?11) z |= 4'b0100; 
	if(x==?20'b1?1?111?1?????00???1) z |= 4'b1000; 
	if(x==?20'b?11?0??10?11????1??1) z |= 4'b0100; 
	if(x==?20'b???1?11?01??00???11?) z |= 4'b0100; 
	if(x==?20'b??1?0??1?1??000??1?1) z |= 4'b0100; 
	if(x==?20'b?????11???01?00111??) z |= 4'b1000; 
	if(x==?20'b?1??1??0??1??000?1?1) z |= 4'b1000; 
	if(x==?20'b?1??0111?110????11??) z |= 4'b1100; 
	if(x==?20'b??1?111???0??000???1) z |= 4'b1000; 
	if(x==?20'b?1?1???1???10?1?111?) z |= 4'b0100; 
	if(x==?20'b111?1?1011???????1??) z |= 4'b1000; 
	if(x==?20'b?11?1???11?0???01??1) z |= 4'b1000; 
	if(x==?20'b??11???1??1?0?1?1?11) z |= 4'b0100; 
	if(x==?20'b?1???1110???000????1) z |= 4'b0100; 
	if(x==?20'b??1?111????0?000???1) z |= 4'b1000; 
	if(x==?20'b1????11???10??00?11?) z |= 4'b1000; 
	if(x==?20'b11??111???00????1?1?) z |= 4'b1000; 
	if(x==?20'b1?1??11?1????1?01??1) z |= 4'b1000; 
	if(x==?20'b?1???111?0??000????1) z |= 4'b0100; 
	if(x==?20'b?1?1?111???100?????1) z |= 4'b0100; 
	if(x==?20'b?????1?011???0?11?11) z |= 4'b1000; 
	if(x==?20'b??11?111???10?0????1) z |= 4'b0100; 
	if(x==?20'b111?11??110?????1???) z |= 4'b1000; 
	if(x==?20'b??11???1??1100??1??1) z |= 4'b0100; 
	if(x==?20'b??11?11100??????1?1?) z |= 4'b0100; 
	if(x==?20'b?1??011???1?0?1?1??1) z |= 4'b0100; 
	if(x==?20'b?11?1??011?????01??1) z |= 4'b1000; 
	if(x==?20'b1?1??1101??0?????11?) z |= 4'b1000; 
	if(x==?20'b?????1??110??000?11?) z |= 4'b1000; 
	if(x==?20'b??1?0?11111??0?????1) z |= 4'b0100; 
	if(x==?20'b1????110?????0001??1) z |= 4'b1000; 
	if(x==?20'b1?1????01????0?0?111) z |= 4'b1000; 
	if(x==?20'b?1??011101????0??11?) z |= 4'b1100; 
	if(x==?20'b??1?1?1011?????0?11?) z |= 4'b1000; 
	if(x==?20'b?11?1?10?1?0?0???1??) z |= 4'b1000; 
	if(x==?20'b????1?10?1???000?11?) z |= 4'b1000; 
	if(x==?20'b???1?1?1??110?0??11?) z |= 4'b0100; 
	if(x==?20'b1????1111?0???0???11) z |= 4'b1000; 
	if(x==?20'b?11????10?110???1??1) z |= 4'b0100; 
	if(x==?20'b?111?1?1??11?1???1??) z |= 4'b0100; 
	if(x==?20'b?1?1011?0??1?????11?) z |= 4'b0100; 
	if(x==?20'b?1??1?101??0?0???11?) z |= 4'b1000; 
	if(x==?20'b??1?1110??10?0???11?) z |= 4'b1100; 
	if(x==?20'b?1??11??110????01?1?) z |= 4'b1000; 
	if(x==?20'b?1??11?0?111??0????1) z |= 4'b1000; 
	if(x==?20'b?11?01?10?1???0??1??) z |= 4'b0100; 
	if(x==?20'b?11101?1??11?????1??) z |= 4'b0100; 
	if(x==?20'b11??1??0??????001?11) z |= 4'b1000; 
	if(x==?20'b?1?10??????10?0??111) z |= 4'b0100; 
	if(x==?20'b???1111??0?1?0????11) z |= 4'b0100; 
	if(x==?20'b????01?1??1?000??11?) z |= 4'b0100; 
	if(x==?20'b??110???1???00??11?1) z |= 4'b0100; 
	if(x==?20'b?11???11011?0???1???) z |= 4'b0100; 
	if(x==?20'b111?1?10???0?????11?) z |= 4'b1000; 
	if(x==?20'b??1?1???0???100?11?1) z |= 4'b0100; 
	if(x==?20'b?11101?10????????11?) z |= 4'b0100; 
	if(x==?20'b?11?11???110???01???) z |= 4'b1000; 
	if(x==?20'b??11???101???00??1?1) z |= 4'b0100; 
	if(x==?20'b?11?0??1??110???1??1) z |= 4'b0100; 
	if(x==?20'b??????1??011000??11?) z |= 4'b0100; 
	if(x==?20'b111??1?0111????????1) z |= 4'b1000; 
	if(x==?20'b?111??11?011????1???) z |= 4'b0100; 
	if(x==?20'b?1?1?11????10?1?1??1) z |= 4'b0100; 
	if(x==?20'b??1?01?10??1??0??11?) z |= 4'b0100; 
	if(x==?20'b???10?11?1???00?1??1) z |= 4'b0100; 
	if(x==?20'b111?11????00????1?1?) z |= 4'b1000; 
	if(x==?20'b??1?1?101????10?11??) z |= 4'b1000; 
	if(x==?20'b?1??01?1??110????11?) z |= 4'b0100; 
	if(x==?20'b11??1?????10?00??1?1) z |= 4'b1000; 
	if(x==?20'b?111??1100??????1?1?) z |= 4'b0100; 
	if(x==?20'b??1???11111?00?????1) z |= 4'b0100; 
	if(x==?20'b11??1???1????0?11?11) z |= 4'b1000; 
	if(x==?20'b1?1??11?1110?????1??) z |= 4'b1000; 
	if(x==?20'b11?????0???1??0011?1) z |= 4'b1000; 
	if(x==?20'b?1110?1??111???????1) z |= 4'b0100; 
	if(x==?20'b1???1?10?????0?0111?) z |= 4'b1000; 
	if(x==?20'b?1??1?1?1??0?0?0?11?) z |= 4'b1000; 
	if(x==?20'b1?1??1101??????0?11?) z |= 4'b1000; 
	if(x==?20'b?1??01?1?0?1?0??11??) z |= 4'b0100; 
	if(x==?20'b?1?1?11?0111?????1??) z |= 4'b0100; 
	if(x==?20'b?11??11??11?11??1???) z |= 4'b0100; 
	if(x==?20'b???101?1????0?0?111?) z |= 4'b0100; 
	if(x==?20'b1?1?111??1???0?0???1) z |= 4'b1000; 
	if(x==?20'b1???111?11?0????1?1?) z |= 4'b1000; 
	if(x==?20'b????011101???0???11?) z |= 4'b0100; 
	if(x==?20'b?1??11???111??00???1) z |= 4'b1000; 
	if(x==?20'b?1?????1???0?00111?1) z |= 4'b1000; 
	if(x==?20'b111?11??11?????01???) z |= 4'b1000; 
	if(x==?20'b111?1???11?0????1??1) z |= 4'b1000; 
	if(x==?20'b?11?0??101???0???1?1) z |= 4'b0100; 
	if(x==?20'b111?11?0???0????1?1?) z |= 4'b1000; 
	if(x==?20'b?1??1?101????0?0?11?) z |= 4'b1000; 
	if(x==?20'b1???111?1?????00??11) z |= 4'b1000; 
	if(x==?20'b1?????101?????00111?) z |= 4'b1000; 
	if(x==?20'b1?1?111????0?00????1) z |= 4'b1000; 
	if(x==?20'b?1?1?1110????00????1) z |= 4'b0100; 
	if(x==?20'b?11??1?1??1?010??1??) z |= 4'b0100; 
	if(x==?20'b????1110??10??0??11?) z |= 4'b1000; 
	if(x==?20'b?1?1011????10????11?) z |= 4'b0100; 
	if(x==?20'b?11?1?1??1???010?1??) z |= 4'b1000; 
	if(x==?20'b??11??11??1?1?0?1?1?) z |= 4'b0100; 
	if(x==?20'b?11????1?001?0??11??) z |= 4'b0100; 
	if(x==?20'b??1??1?10??10?0??11?) z |= 4'b0100; 
	if(x==?20'b11??1110?11?????1???) z |= 4'b1000; 
	if(x==?20'b?11?0??1????0?1?1?11) z |= 4'b0100; 
	if(x==?20'b?11?1??0??10??0??1?1) z |= 4'b1000; 
	if(x==?20'b?1?1?111??1?0?0????1) z |= 4'b0100; 
	if(x==?20'b111?1??011??????1??1) z |= 4'b1000; 
	if(x==?20'b?????11?110??10?11??) z |= 4'b1000; 
	if(x==?20'b11???11?1110????1???) z |= 4'b1000; 
	if(x==?20'b11??11???1???0?11?1?) z |= 4'b1000; 
	if(x==?20'b?1?????10??1?10??111) z |= 4'b0100; 
	if(x==?20'b?????11011????001??1) z |= 4'b1000; 
	if(x==?20'b??110111?11?????1???) z |= 4'b0100; 
	if(x==?20'b?1???1111?0????0??11) z |= 4'b1000; 
	if(x==?20'b1?1??11??1???1?01??1) z |= 4'b1000; 
	if(x==?20'b????111??0??000???11) z |= 4'b0100; 
	if(x==?20'b?????111??0??000??11) z |= 4'b1000; 
	if(x==?20'b1?1?1?1011???????11?) z |= 4'b1000; 
	if(x==?20'b??1?1???1??0?01??111) z |= 4'b1000; 
	if(x==?20'b???101?????100??111?) z |= 4'b0100; 
	if(x==?20'b?1??0?11011?????1?1?) z |= 4'b0100; 
	if(x==?20'b???1?1110?11????1?1?) z |= 4'b0100; 
	if(x==?20'b??1???11??110?1?1?1?) z |= 4'b0100; 
	if(x==?20'b??1?11?0?110????1?1?) z |= 4'b1000; 
	if(x==?20'b???1?111???100????11) z |= 4'b0100; 
	if(x==?20'b??1?01?1???1?01?11??) z |= 4'b0100; 
	if(x==?20'b11???1101??????01?1?) z |= 4'b1000; 
	if(x==?20'b?111???10?11????1??1) z |= 4'b0100; 
	if(x==?20'b??11?11?0111????1???) z |= 4'b0100; 
	if(x==?20'b?111??11??110???1???) z |= 4'b0100; 
	if(x==?20'b?1?1???1????010?111?) z |= 4'b0100; 
	if(x==?20'b??1?01?1???10?0??11?) z |= 4'b0100; 
	if(x==?20'b??1?111??0?10?????11) z |= 4'b0100; 
	if(x==?20'b??1?1?0???0??00?111?) z |= 4'b1000; 
	if(x==?20'b????11?0111???0???11) z |= 4'b1000; 
	if(x==?20'b111???1???00??0???11) z |= 4'b1000; 
	if(x==?20'b?111?1??00???0????11) z |= 4'b0100; 
	if(x==?20'b?11??11??11???111???) z |= 4'b1000; 
	if(x==?20'b?11????101??00???1?1) z |= 4'b0100; 
	if(x==?20'b11??????11???000?1?1) z |= 4'b1000; 
	if(x==?20'b??11011????10???1?1?) z |= 4'b0100; 
	if(x==?20'b?111??11011?????1???) z |= 4'b0100; 
	if(x==?20'b1?1?11??11?0????1?1?) z |= 4'b1000; 
	if(x==?20'b1?1?1????????010111?) z |= 4'b1000; 
	if(x==?20'b111?11???110????1???) z |= 4'b1000; 
	if(x==?20'b1????1??11???0?11?11) z |= 4'b1000; 
	if(x==?20'b?1??0?11?1??00??1??1) z |= 4'b0100; 
	if(x==?20'b?1110??1??11????1??1) z |= 4'b0100; 
	if(x==?20'b?1???0?1?0???00?111?) z |= 4'b0100; 
	if(x==?20'b?11?01101??1?????11?) z |= 4'b1100; 
	if(x==?20'b?11?1?????10??00?1?1) z |= 4'b1000; 
	if(x==?20'b?1?1?11???1?0?1?1??1) z |= 4'b0100; 
	if(x==?20'b??1?11?0???0?00?1??1) z |= 4'b1000; 
	if(x==?20'b????0?11?111?0????11) z |= 4'b0100; 
	if(x==?20'b?1?101?1??11?????11?) z |= 4'b0100; 
	if(x==?20'b1?1?1???1????0?1111?) z |= 4'b1000; 
	if(x==?20'b1?1?11?011??????1?1?) z |= 4'b1000; 
	if(x==?20'b??11??11111??0?????1) z |= 4'b0100; 
	if(x==?20'b1?1?111??????000???1) z |= 4'b1000; 
	if(x==?20'b1?1?1?1?11?????0?11?) z |= 4'b1000; 
	if(x==?20'b1???1?1??1???000?11?) z |= 4'b1000; 
	if(x==?20'b11???110?1?0????1?1?) z |= 4'b1000; 
	if(x==?20'b1?1?1????10??00?11??) z |= 4'b1000; 
	if(x==?20'b??11011?0?1?????1?1?) z |= 4'b0100; 
	if(x==?20'b?1?1?111????000????1) z |= 4'b0100; 
	if(x==?20'b?1?1??110?11????1?1?) z |= 4'b0100; 
	if(x==?20'b??11??????11000??1?1) z |= 4'b0100; 
	if(x==?20'b11???1?0111???????11) z |= 4'b1000; 
	if(x==?20'b11??1?1?1??0?0???11?) z |= 4'b1000; 
	if(x==?20'b??1?11??00???00?1?11) z |= 4'b1100; 
	if(x==?20'b1?1?1?1?1??0??0??11?) z |= 4'b1000; 
	if(x==?20'b1????1?1?1???000?11?) z |= 4'b1000; 
	if(x==?20'b?????11??011?01?11??) z |= 4'b0100; 
	if(x==?20'b11??1????1???0?11?11) z |= 4'b1000; 
	if(x==?20'b11??11???111??0????1) z |= 4'b1000; 
	if(x==?20'b?1????11??00?00?1?11) z |= 4'b1100; 
	if(x==?20'b?111?1??1???0?1?11??) z |= 4'b0100; 
	if(x==?20'b????11??111???00??11) z |= 4'b1000; 
	if(x==?20'b11??1????1?0?00?11??) z |= 4'b1000; 
	if(x==?20'b??110?11?1?1????1?1?) z |= 4'b0100; 
	if(x==?20'b111?111?1?0???????1?) z |= 4'b1000; 
	if(x==?20'b?????1101????0001??1) z |= 4'b1000; 
	if(x==?20'b???1?1?1??1?000??11?) z |= 4'b0100; 
	if(x==?20'b??1????1??110?1?1?11) z |= 4'b0100; 
	if(x==?20'b??110?1??111??????11) z |= 4'b0100; 
	if(x==?20'b11??1?101????0???11?) z |= 4'b1000; 
	if(x==?20'b1?1?1?101?????0??11?) z |= 4'b1000; 
	if(x==?20'b?1110????0?1????1?11) z |= 4'b0100; 
	if(x==?20'b??11???10?1??00?11??) z |= 4'b0100; 
	if(x==?20'b?1?1011?0?????0??11?) z |= 4'b0100; 
	if(x==?20'b?1?10?11??11????1?1?) z |= 4'b0100; 
	if(x==?20'b?1?1???1?01??00?11??) z |= 4'b0100; 
	if(x==?20'b?1?1?1?10??1?0???11?) z |= 4'b0100; 
	if(x==?20'b111???1????1??1011??) z |= 4'b1000; 
	if(x==?20'b1?1??110???0?0???11?) z |= 4'b1000; 
	if(x==?20'b??11?1?10??1??0??11?) z |= 4'b0100; 
	if(x==?20'b111?111?1??0??????1?) z |= 4'b1000; 
	if(x==?20'b?111??1?0???00????11) z |= 4'b0100; 
	if(x==?20'b??1?1?10?1???0?0?11?) z |= 4'b1000; 
	if(x==?20'b??????11?11100????11) z |= 4'b0100; 
	if(x==?20'b????011????1000?1??1) z |= 4'b0100; 
	if(x==?20'b?1?1?1?1??110????11?) z |= 4'b0100; 
	if(x==?20'b?11???1?011?0?0??1??) z |= 4'b0100; 
	if(x==?20'b1????111??0??00???11) z |= 4'b1000; 
	if(x==?20'b???1111??0???00???11) z |= 4'b0100; 
	if(x==?20'b?11?01??1???10??11??) z |= 4'b0100; 
	if(x==?20'b??1?0?1?011??0??1??1) z |= 4'b0100; 
	if(x==?20'b111?1????????1?01?11) z |= 4'b1000; 
	if(x==?20'b1????11?1110????11??) z |= 4'b1000; 
	if(x==?20'b?11????1001???0?11??) z |= 4'b0100; 
	if(x==?20'b?11?1?101??0?????11?) z |= 4'b1000; 
	if(x==?20'b11???11??1?0???01?1?) z |= 4'b1000; 
	if(x==?20'b11??1?101????0??11??) z |= 4'b1000; 
	if(x==?20'b?11??1???110?0?0?1??) z |= 4'b1000; 
	if(x==?20'b??11?11?0?1?0???1?1?) z |= 4'b0100; 
	if(x==?20'b111??1?????0??00??11) z |= 4'b1000; 
	if(x==?20'b?1?101?1???1?0???11?) z |= 4'b0100; 
	if(x==?20'b?111?1110??1??????1?) z |= 4'b0100; 
	if(x==?20'b?111?111?0?1??????1?) z |= 4'b0100; 
	if(x==?20'b??1101?1???1??0??11?) z |= 4'b0100; 
	if(x==?20'b?1???1?0?110??0?1??1) z |= 4'b1000; 
	if(x==?20'b1?1?1??011??????1?11) z |= 4'b1000; 
	if(x==?20'b???1?11?0111????11??) z |= 4'b0100; 
	if(x==?20'b?1??111?00????0???11) z |= 4'b0100; 
	if(x==?20'b?1110?1?????00????11) z |= 4'b0100; 
	if(x==?20'b?11?11??1?00????1?1?) z |= 4'b1000; 
	if(x==?20'b?1??01?1??1?0?0??11?) z |= 4'b0100; 
	if(x==?20'b??1??111??00?0????11) z |= 4'b1000; 
	if(x==?20'b11???110?1?????01?1?) z |= 4'b1000; 
	if(x==?20'b?111???101???0???1?1) z |= 4'b0100; 
	if(x==?20'b????1111????111????1) z |= 4'b0100; 
	if(x==?20'b111??1?0??????00??11) z |= 4'b1000; 
	if(x==?20'b11??1?1?1????0?0?11?) z |= 4'b1000; 
	if(x==?20'b????1?101????0?0111?) z |= 4'b1000; 
	if(x==?20'b?11?01?10??1?????11?) z |= 4'b0100; 
	if(x==?20'b11????1?11?0?0??1??1) z |= 4'b1000; 
	if(x==?20'b??11011???1?0???1?1?) z |= 4'b0100; 
	if(x==?20'b11????1?11?0??0?1??1) z |= 4'b1000; 
	if(x==?20'b????1?1101???00??11?) z |= 4'b0100; 
	if(x==?20'b?111???1????0?1?1?11) z |= 4'b0100; 
	if(x==?20'b111?1?????10??0??1?1) z |= 4'b1000; 
	if(x==?20'b????0?11?1?1?00?1??1) z |= 4'b0100; 
	if(x==?20'b??????101??0?00??111) z |= 4'b1000; 
	if(x==?20'b??1?111?11???0?0???1) z |= 4'b1000; 
	if(x==?20'b?11???1100?1????1?1?) z |= 4'b0100; 
	if(x==?20'b1????11?11????001??1) z |= 4'b1000; 
	if(x==?20'b111??1??11???0?0?1??) z |= 4'b1000; 
	if(x==?20'b?11???10???1??0111??) z |= 4'b1000; 
	if(x==?20'b1?1?1?10???????0111?) z |= 4'b1000; 
	if(x==?20'b??1???1?011?00??1??1) z |= 4'b0100; 
	if(x==?20'b?11?11?01??0????1?1?) z |= 4'b1000; 
	if(x==?20'b????1111?????111???1) z |= 4'b1000; 
	if(x==?20'b?1?1??11011?????1?1?) z |= 4'b0100; 
	if(x==?20'b?11?1?1?1??0???0?11?) z |= 4'b1000; 
	if(x==?20'b1?1?11???110????1?1?) z |= 4'b1000; 
	if(x==?20'b??1?111?1??0?00????1) z |= 4'b1000; 
	if(x==?20'b?1?10??1??11????1?11) z |= 4'b0100; 
	if(x==?20'b?1?101?1????0???111?) z |= 4'b0100; 
	if(x==?20'b????11?1??10?00??11?) z |= 4'b1000; 
	if(x==?20'b??11?1??0?11?0??1??1) z |= 4'b0100; 
	if(x==?20'b????01??0??1?00??111) z |= 4'b0100; 
	if(x==?20'b111?1??0?1????0???11) z |= 4'b1000; 
	if(x==?20'b111?111?111?????????) z |= 4'b1000; 
	if(x==?20'b??11?1??0?11??0?1??1) z |= 4'b0100; 
	if(x==?20'b??11?1?1???10?0??11?) z |= 4'b0100; 
	if(x==?20'b????01?1???10?0?111?) z |= 4'b0100; 
	if(x==?20'b?1???1???110??001??1) z |= 4'b1000; 
	if(x==?20'b?11?1????1?0??0011??) z |= 4'b1000; 
	if(x==?20'b1???11??111???0???11) z |= 4'b1000; 
	if(x==?20'b11????101??????0111?) z |= 4'b1000; 
	if(x==?20'b?????11??1?0?0001??1) z |= 4'b1000; 
	if(x==?20'b?1??11??11???0?11?1?) z |= 4'b1000; 
	if(x==?20'b?11?1?101??????0?11?) z |= 4'b1000; 
	if(x==?20'b1???111??????000??11) z |= 4'b1000; 
	if(x==?20'b?11????10?1?00??11??) z |= 4'b0100; 
	if(x==?20'b?1??1?10?????000?11?) z |= 4'b1000; 
	if(x==?20'b?????11?0?1?000?1??1) z |= 4'b0100; 
	if(x==?20'b?1110??1??1??0????11) z |= 4'b0100; 
	if(x==?20'b?111??1???110?0??1??) z |= 4'b0100; 
	if(x==?20'b?1???1110??1?00????1) z |= 4'b0100; 
	if(x==?20'b?11??1?10??10????11?) z |= 4'b0100; 
	if(x==?20'b?????1?011????001?11) z |= 4'b1000; 
	if(x==?20'b???1?111????000???11) z |= 4'b0100; 
	if(x==?20'b??1?01?1????000??11?) z |= 4'b0100; 
	if(x==?20'b??1?111?0???00????11) z |= 4'b0100; 
	if(x==?20'b?11?1??0?????0?11?11) z |= 4'b1000; 
	if(x==?20'b?1???111??110?0????1) z |= 4'b0100; 
	if(x==?20'b?????110?1???0001??1) z |= 4'b1000; 
	if(x==?20'b?1??111??0??00????11) z |= 4'b0100; 
	if(x==?20'b?1???111??0??0?0??11) z |= 4'b1000; 
	if(x==?20'b1?1?1?10?1???0???11?) z |= 4'b1000; 
	if(x==?20'b??1?111??0??0?0???11) z |= 4'b0100; 
	if(x==?20'b??1??1111110????11??) z |= 4'b1100; 
	if(x==?20'b??1??111??0???00??11) z |= 4'b1000; 
	if(x==?20'b???1??11?111?0????11) z |= 4'b0100; 
	if(x==?20'b?111?111?111????????) z |= 4'b0100; 
	if(x==?20'b??????1?1??0?000?111) z |= 4'b1000; 
	if(x==?20'b???1011????1?00?1??1) z |= 4'b0100; 
	if(x==?20'b??1101?????10???111?) z |= 4'b0100; 
	if(x==?20'b??1?111????0?0?0??11) z |= 4'b1000; 
	if(x==?20'b?1??111?0111????11??) z |= 4'b1100; 
	if(x==?20'b?11?1?101??????011??) z |= 4'b1000; 
	if(x==?20'b?1???1110???0?0???11) z |= 4'b0100; 
	if(x==?20'b????011???1?000?1??1) z |= 4'b0100; 
	if(x==?20'b?11?1?101??1?0???11?) z |= 4'b1100; 
	if(x==?20'b?11?01?1???10????11?) z |= 4'b0100; 
	if(x==?20'b?11?11??1110????1???) z |= 4'b1000; 
	if(x==?20'b?1???111???0??00??11) z |= 4'b1000; 
	if(x==?20'b11??11???10???0?1?1?) z |= 4'b1000; 
	if(x==?20'b??1?11?0111???????11) z |= 4'b1000; 
	if(x==?20'b?????1??0??1000??111) z |= 4'b0100; 
	if(x==?20'b111?1????1????00??11) z |= 4'b1000; 
	if(x==?20'b????11?1?1???000?11?) z |= 4'b1000; 
	if(x==?20'b??1??1111??0?00???11) z |= 4'b1100; 
	if(x==?20'b?11?01?11??1??0??11?) z |= 4'b1100; 
	if(x==?20'b?1?101?1??1???0??11?) z |= 4'b0100; 
	if(x==?20'b?1??111?0??1?00???11) z |= 4'b1100; 
	if(x==?20'b1????11?1????0001??1) z |= 4'b1000; 
	if(x==?20'b?11?011?011?????1???) z |= 4'b0100; 
	if(x==?20'b??1?111?1????000???1) z |= 4'b1000; 
	if(x==?20'b?11???110111????1???) z |= 4'b0100; 
	if(x==?20'b?11???1?11?0???01??1) z |= 4'b1000; 
	if(x==?20'b????1?1?11???000?11?) z |= 4'b1000; 
	if(x==?20'b1???1?101????0??111?) z |= 4'b1000; 
	if(x==?20'b?111???1??1?00????11) z |= 4'b0100; 
	if(x==?20'b?1???11011?0????1?1?) z |= 4'b1000; 
	if(x==?20'b?????11?01??000??11?) z |= 4'b0100; 
	if(x==?20'b??11??11?01??0??1?1?) z |= 4'b0100; 
	if(x==?20'b?11??110?110????1???) z |= 4'b1000; 
	if(x==?20'b?11?01?1???10???11??) z |= 4'b0100; 
	if(x==?20'b111?11??111????????1) z |= 4'b1000; 
	if(x==?20'b?1??0?11?111??????11) z |= 4'b0100; 
	if(x==?20'b?1???11???110?1?1??1) z |= 4'b0100; 
	if(x==?20'b111?111??????0?0???1) z |= 4'b1000; 
	if(x==?20'b?1??1???11???0?11?11) z |= 4'b1000; 
	if(x==?20'b11??1?1111??????1??1) z |= 4'b1000; 
	if(x==?20'b1?1?1?1??1???0?0?11?) z |= 4'b1000; 
	if(x==?20'b???1?11????1000?1??1) z |= 4'b0100; 
	if(x==?20'b11??1???1?????001?11) z |= 4'b1000; 
	if(x==?20'b?????11???10?000?11?) z |= 4'b1000; 
	if(x==?20'b?111?111????0?0????1) z |= 4'b0100; 
	if(x==?20'b111?1?1?1??0?????11?) z |= 4'b1000; 
	if(x==?20'b??1?011?0?11????1?1?) z |= 4'b0100; 
	if(x==?20'b?11??1??0?110???1??1) z |= 4'b0100; 
	if(x==?20'b?1???111???1000????1) z |= 4'b0100; 
	if(x==?20'b11???10??10????0?1??) z |= 4'b1000; 
	if(x==?20'b?11?11??110??0??1???) z |= 4'b1000; 
	if(x==?20'b?11?11??110???0?1???) z |= 4'b1000; 
	if(x==?20'b?11?1?1?11???01??1??) z |= 4'b1000; 
	if(x==?20'b?111??11?111???????1) z |= 4'b0100; 
	if(x==?20'b???101?1???1??0?111?) z |= 4'b0100; 
	if(x==?20'b?1?1?1?1??1?0?0??11?) z |= 4'b0100; 
	if(x==?20'b??11?01??01?0????1??) z |= 4'b0100; 
	if(x==?20'b111?1?101????????11?) z |= 4'b1000; 
	if(x==?20'b111??11011??????1???) z |= 4'b1000; 
	if(x==?20'b?????1?1??11000??11?) z |= 4'b0100; 
	if(x==?20'b?????1111?0??00???11) z |= 4'b1000; 
	if(x==?20'b?111?1?10??1?????11?) z |= 4'b0100; 
	if(x==?20'b?1???11?11?0???01?1?) z |= 4'b1000; 
	if(x==?20'b?????????111111???11) z |= 4'b0100; 
	if(x==?20'b??1111?1??11????1??1) z |= 4'b0100; 
	if(x==?20'b?11??1?1??11?10??1??) z |= 4'b0100; 
	if(x==?20'b????????111??111??11) z |= 4'b1000; 
	if(x==?20'b11??111?111???????1?) z |= 4'b1000; 
	if(x==?20'b1?1??1101??1????11??) z |= 4'b1000; 
	if(x==?20'b?1?1011?1??1????11??) z |= 4'b0100; 
	if(x==?20'b??11111?0????0????11) z |= 4'b0100; 
	if(x==?20'b11???111??0??0????11) z |= 4'b1000; 
	if(x==?20'b?1?1111??0???0????11) z |= 4'b0100; 
	if(x==?20'b1?1??111??0???0???11) z |= 4'b1000; 
	if(x==?20'b??11111??0????0???11) z |= 4'b0100; 
	if(x==?20'b1?????1?1??0?00??111) z |= 4'b1000; 
	if(x==?20'b??11??11?1??00??1?1?) z |= 4'b0100; 
	if(x==?20'b111???1????1?0?111??) z |= 4'b1000; 
	if(x==?20'b????111??0?1?00???11) z |= 4'b0100; 
	if(x==?20'b?1???11011?????01?1?) z |= 4'b1000; 
	if(x==?20'b??1?0???1???000?11?1) z |= 4'b0100; 
	if(x==?20'b111?1?101???????11??) z |= 4'b1000; 
	if(x==?20'b???1011???1??00?1??1) z |= 4'b0100; 
	if(x==?20'b??1??11?0?110???1?1?) z |= 4'b0100; 
	if(x==?20'b?11???11?011?0??1???) z |= 4'b0100; 
	if(x==?20'b11??11????1???001?1?) z |= 4'b1000; 
	if(x==?20'b????11111?1??00?1??1) z |= 4'b1100; 
	if(x==?20'b?11101?1???1?????11?) z |= 4'b0100; 
	if(x==?20'b?111011???11????1???) z |= 4'b0100; 
	if(x==?20'b11???111???0??0???11) z |= 4'b1000; 
	if(x==?20'b?11???11?011??0?1???) z |= 4'b0100; 
	if(x==?20'b?1??011?0??1??0?11??) z |= 4'b0100; 
	if(x==?20'b?1?1???1???1?10?111?) z |= 4'b0100; 
	if(x==?20'b???1?1??0??1?00??111) z |= 4'b0100; 
	if(x==?20'b?11?11????00?0??1?1?) z |= 4'b1000; 
	if(x==?20'b?11?11????00??0?1?1?) z |= 4'b1000; 
	if(x==?20'b?11?1??11????10?11??) z |= 4'b1000; 
	if(x==?20'b????1111?1?1?00?1??1) z |= 4'b1100; 
	if(x==?20'b?11???1100???0??1?1?) z |= 4'b0100; 
	if(x==?20'b??1?01???1??000??11?) z |= 4'b0100; 
	if(x==?20'b??11?111?111??????1?) z |= 4'b0100; 
	if(x==?20'b?11???1100????0?1?1?) z |= 4'b0100; 
	if(x==?20'b11??1???11???00?1??1) z |= 4'b1000; 
	if(x==?20'b?11?11???1???1?01?1?) z |= 4'b1000; 
	if(x==?20'b?1?????0???1?00011?1) z |= 4'b1000; 
	if(x==?20'b??1?1?101??????0111?) z |= 4'b1000; 
	if(x==?20'b1?1?111?1????00????1) z |= 4'b1000; 
	if(x==?20'b11??1?1??????000?11?) z |= 4'b1000; 
	if(x==?20'b111???1?11?0????1??1) z |= 4'b1000; 
	if(x==?20'b?1????10??1??000?11?) z |= 4'b1000; 
	if(x==?20'b??1??1101????01?11??) z |= 4'b1000; 
	if(x==?20'b1?1?11???????000?11?) z |= 4'b1000; 
	if(x==?20'b?1??1?1101???0???11?) z |= 4'b0100; 
	if(x==?20'b1????1??11????001?11) z |= 4'b1000; 
	if(x==?20'b??1?011???110???1?1?) z |= 4'b0100; 
	if(x==?20'b???1?11?01???00??11?) z |= 4'b0100; 
	if(x==?20'b?1?1??11????000??11?) z |= 4'b0100; 
	if(x==?20'b?11101?1???1????11??) z |= 4'b0100; 
	if(x==?20'b??11?1?1????000??11?) z |= 4'b0100; 
	if(x==?20'b?11????1???10?1?1?11) z |= 4'b0100; 
	if(x==?20'b111?1?1???0???0???11) z |= 4'b1000; 
	if(x==?20'b?11?1???11?0?0??1??1) z |= 4'b1000; 
	if(x==?20'b?11?1???11?0??0?1??1) z |= 4'b1000; 
	if(x==?20'b?11?1?1????0?0?0?11?) z |= 4'b1000; 
	if(x==?20'b????111?1????000??11) z |= 4'b1000; 
	if(x==?20'b1????11???10?00??11?) z |= 4'b1000; 
	if(x==?20'b1?1??1??1????000?11?) z |= 4'b1000; 
	if(x==?20'b1?1?111???10????11??) z |= 4'b1000; 
	if(x==?20'b??1?11?1??10??0??11?) z |= 4'b1000; 
	if(x==?20'b?11??1?10???0?0??11?) z |= 4'b0100; 
	if(x==?20'b?111?1??0?11????1??1) z |= 4'b0100; 
	if(x==?20'b?1?1?111???1?00????1) z |= 4'b0100; 
	if(x==?20'b?1??01?1???10???111?) z |= 4'b0100; 
	if(x==?20'b????????111?111???1?) z |= 4'b0010; 
	if(x==?20'b?111?1?1?0???0????11) z |= 4'b0100; 
	if(x==?20'b1?1?11??111???????11) z |= 4'b1000; 
	if(x==?20'b?11?1??011???0??1??1) z |= 4'b1000; 
	if(x==?20'b??11???1??11?00?1??1) z |= 4'b0100; 
	if(x==?20'b11??1????1????001?11) z |= 4'b1000; 
	if(x==?20'b?11?1??011????0?1??1) z |= 4'b1000; 
	if(x==?20'b11??111??????0?0??11) z |= 4'b1000; 
	if(x==?20'b1?1?111???????00??11) z |= 4'b1000; 
	if(x==?20'b1?1???10??????00111?) z |= 4'b1000; 
	if(x==?20'b?1?101??????00??111?) z |= 4'b0100; 
	if(x==?20'b?11???11??1?0?1?1?1?) z |= 4'b0100; 
	if(x==?20'b?1?1??1????1000??11?) z |= 4'b0100; 
	if(x==?20'b11??11???????0001?1?) z |= 4'b1000; 
	if(x==?20'b?1?1?111????00????11) z |= 4'b0100; 
	if(x==?20'b?111?11?011?????1???) z |= 4'b0100; 
	if(x==?20'b??11??11????000?1?1?) z |= 4'b0100; 
	if(x==?20'b1?1??11?1?10????11??) z |= 4'b1000; 
	if(x==?20'b??11?111????0?0???11) z |= 4'b0100; 
	if(x==?20'b?11????10?11?0??1??1) z |= 4'b0100; 
	if(x==?20'b11???11?11?0????1?1?) z |= 4'b1000; 
	if(x==?20'b?????111???1000???11) z |= 4'b0100; 
	if(x==?20'b?11????10?11??0?1??1) z |= 4'b0100; 
	if(x==?20'b111??11??110????1???) z |= 4'b1000; 
	if(x==?20'b?11?111??0??0?????11) z |= 4'b0100; 
	if(x==?20'b?11??111??0????0??11) z |= 4'b1000; 
	if(x==?20'b?1??11??110???0?1?1?) z |= 4'b1000; 
	if(x==?20'b?1?1??11?111??????11) z |= 4'b0100; 
	if(x==?20'b??1???1?1??0??00?111) z |= 4'b1000; 
	if(x==?20'b?11????1???0?10?11?1) z |= 4'b1000; 
	if(x==?20'b11???11011??????1?1?) z |= 4'b1000; 
	if(x==?20'b?11???11011??0??1???) z |= 4'b0100; 
	if(x==?20'b??110??1?????00?1?11) z |= 4'b0100; 
	if(x==?20'b??110???1????00?11?1) z |= 4'b0100; 
	if(x==?20'b?11?11???110?0??1???) z |= 4'b1000; 
	if(x==?20'b?11???11011???0?1???) z |= 4'b0100; 
	if(x==?20'b111??1?01?????0???11) z |= 4'b1000; 
	if(x==?20'b?1???1??0??100???111) z |= 4'b0100; 
	if(x==?20'b?11?0??1??11?0??1??1) z |= 4'b0100; 
	if(x==?20'b?11?11???110??0?1???) z |= 4'b1000; 
	if(x==?20'b??11?11?0?11????1?1?) z |= 4'b0100; 
	if(x==?20'b?1??011?1?1??00?1??1) z |= 4'b1100; 
	if(x==?20'b??1??1101?1??00?1??1) z |= 4'b1100; 
	if(x==?20'b?11?0??1??11??0?1??1) z |= 4'b0100; 
	if(x==?20'b?????????111?111??1?) z |= 4'b0001; 
	if(x==?20'b?11?1???0????01?11?1) z |= 4'b0100; 
	if(x==?20'b?11??1111??0?0????11) z |= 4'b1100; 
	if(x==?20'b??1??11?11???0?11??1) z |= 4'b1000; 
	if(x==?20'b111?1?10?1??????11??) z |= 4'b1000; 
	if(x==?20'b?1??011??1?1?00?1??1) z |= 4'b1100; 
	if(x==?20'b?11?1???11????001??1) z |= 4'b1000; 
	if(x==?20'b?1110?1????1?0????11) z |= 4'b0100; 
	if(x==?20'b??1??110?1?1?00?1??1) z |= 4'b1100; 
	if(x==?20'b?11?111?1????0?0???1) z |= 4'b1000; 
	if(x==?20'b?11?111?0??1??0???11) z |= 4'b1100; 
	if(x==?20'b???1?11???1?000??11?) z |= 4'b0100; 
	if(x==?20'b??1?1?1?11???0?0?11?) z |= 4'b1000; 
	if(x==?20'b?1????1???110?1?1?11) z |= 4'b0100; 
	if(x==?20'b11?????0???1?00?11?1) z |= 4'b1000; 
	if(x==?20'b??1???11111??00????1) z |= 4'b0100; 
	if(x==?20'b?1???11?01??00???11?) z |= 4'b0100; 
	if(x==?20'b1?1?1?101???????111?) z |= 4'b1000; 
	if(x==?20'b111?11???????0?0??11) z |= 4'b1000; 
	if(x==?20'b??1???11?011?0??1?1?) z |= 4'b0100; 
	if(x==?20'b??11011???11????1?1?) z |= 4'b0100; 
	if(x==?20'b?1???1?0111???0???11) z |= 4'b1000; 
	if(x==?20'b1?1??1101????0???11?) z |= 4'b1000; 
	if(x==?20'b??1???11?011??0?1?1?) z |= 4'b0100; 
	if(x==?20'b?111??11????0?0???11) z |= 4'b0100; 
	if(x==?20'b111????01??1????1?11) z |= 4'b1000; 
	if(x==?20'b?1???10?110????0?1??) z |= 4'b1000; 
	if(x==?20'b1?1??1101?????0??11?) z |= 4'b1000; 
	if(x==?20'b?1??11???111?00????1) z |= 4'b1000; 
	if(x==?20'b?1110?11?1??????1?1?) z |= 4'b0100; 
	if(x==?20'b?11101?1??1?????11??) z |= 4'b0100; 
	if(x==?20'b111?11??11???0??1???) z |= 4'b1000; 
	if(x==?20'b?1???1??1110??0?1??1) z |= 4'b1000; 
	if(x==?20'b11??1????????0001?11) z |= 4'b1000; 
	if(x==?20'b?11????1??1?0?1?1?11) z |= 4'b0100; 
	if(x==?20'b111?11??11????0?1???) z |= 4'b1000; 
	if(x==?20'b??1??11???10??00?11?) z |= 4'b1000; 
	if(x==?20'b?11?111???00????1?1?) z |= 4'b1000; 
	if(x==?20'b??1?0?1??111?0????11) z |= 4'b0100; 
	if(x==?20'b11???11?11?????01?1?) z |= 4'b1000; 
	if(x==?20'b??1???1?0111?0??1??1) z |= 4'b0100; 
	if(x==?20'b1???111?1????00???11) z |= 4'b1000; 
	if(x==?20'b1?????101????00?111?) z |= 4'b1000; 
	if(x==?20'b??11???1????000?1?11) z |= 4'b0100; 
	if(x==?20'b??11????1???000?11?1) z |= 4'b0100; 
	if(x==?20'b?11??111???10?0????1) z |= 4'b0100; 
	if(x==?20'b111??1??1?????00??11) z |= 4'b1000; 
	if(x==?20'b?11????1??1100??1??1) z |= 4'b0100; 
	if(x==?20'b?11??11100??????1?1?) z |= 4'b0100; 
	if(x==?20'b?1?1011????1?0???11?) z |= 4'b0100; 
	if(x==?20'b111??1??111???0????1) z |= 4'b1000; 
	if(x==?20'b?1?101?1???1????111?) z |= 4'b0100; 
	if(x==?20'b?1?1011????1??0??11?) z |= 4'b0100; 
	if(x==?20'b?1??011?????000?1??1) z |= 4'b0100; 
	if(x==?20'b??1??110?????0001??1) z |= 4'b1000; 
	if(x==?20'b?1???1111?0??0????11) z |= 4'b1000; 
	if(x==?20'b?111??1????100????11) z |= 4'b0100; 
	if(x==?20'b??1??1111?0???0???11) z |= 4'b1000; 
	if(x==?20'b?1???1?1??110?0??11?) z |= 4'b0100; 
	if(x==?20'b??1??01??0110????1??) z |= 4'b0100; 
	if(x==?20'b?1??11??11????001?1?) z |= 4'b1000; 
	if(x==?20'b11?????????1?00011?1) z |= 4'b1000; 
	if(x==?20'b?111??1??111?0?????1) z |= 4'b0100; 
	if(x==?20'b???101?????1?00?111?) z |= 4'b0100; 
	if(x==?20'b11???1101????0??1?1?) z |= 4'b1000; 
	if(x==?20'b11???1101?????0?1?1?) z |= 4'b1000; 
	if(x==?20'b???1?111???1?00???11) z |= 4'b0100; 
	if(x==?20'b?111??11??11?0??1???) z |= 4'b0100; 
	if(x==?20'b??11?11???110???1?1?) z |= 4'b0100; 
	if(x==?20'b?1???1??111???00??11) z |= 4'b1000; 
	if(x==?20'b?111??11??11??0?1???) z |= 4'b0100; 
	if(x==?20'b?1???1111??0??0???11) z |= 4'b1000; 
	if(x==?20'b?11?1??0??????001?11) z |= 4'b1000; 
	if(x==?20'b??1?111?0??1?0????11) z |= 4'b0100; 
	if(x==?20'b111?1???11????0???11) z |= 4'b1000; 
	if(x==?20'b?1??111??0?1?0????11) z |= 4'b0100; 
	if(x==?20'b?11?0???1???00??11?1) z |= 4'b0100; 
	if(x==?20'b??1?111??0?1??0???11) z |= 4'b0100; 
	if(x==?20'b??1???1??11100????11) z |= 4'b0100; 
	if(x==?20'b??11011????1?0??1?1?) z |= 4'b0100; 
	if(x==?20'b?11????101???00??1?1) z |= 4'b0100; 
	if(x==?20'b????011???11?00?1??1) z |= 4'b0100; 
	if(x==?20'b??11011????1??0?1?1?) z |= 4'b0100; 
	if(x==?20'b?1??1?1?1????000?11?) z |= 4'b1000; 
	if(x==?20'b?1??0?11?1???00?1??1) z |= 4'b0100; 
	if(x==?20'b?11?1?????10?00??1?1) z |= 4'b1000; 
	if(x==?20'b?111?1??1????10?11??) z |= 4'b0100; 
	if(x==?20'b?????11?11???0001??1) z |= 4'b1000; 
	if(x==?20'b?11????0???1??0011?1) z |= 4'b1000; 
	if(x==?20'b??1?1?10?????0?0111?) z |= 4'b1000; 
	if(x==?20'b1?1?1?1?11???0???11?) z |= 4'b1000; 
	if(x==?20'b?????1?1001?1???11??) z |= 4'b0100; 
	if(x==?20'b?111???1??11?0????11) z |= 4'b0100; 
	if(x==?20'b????1?1??100???111??) z |= 4'b1000; 
	if(x==?20'b??1?111?11?0????1?1?) z |= 4'b1000; 
	if(x==?20'b?1??01?1????0?0?111?) z |= 4'b0100; 
	if(x==?20'b??1??1?1???1000??11?) z |= 4'b0100; 
	if(x==?20'b????11??111??00???11) z |= 4'b1000; 
	if(x==?20'b?1??1???11????001?11) z |= 4'b1000; 
	if(x==?20'b?1??111?1????0?0??11) z |= 4'b1000; 
	if(x==?20'b?1????101????0?0111?) z |= 4'b1000; 
	if(x==?20'b??1?111?1?????00??11) z |= 4'b1000; 
	if(x==?20'b??1???101?????00111?) z |= 4'b1000; 
	if(x==?20'b?????11???11000?1??1) z |= 4'b0100; 
	if(x==?20'b1?1??110?????00?1??1) z |= 4'b1000; 
	if(x==?20'b?1?1011??????00?1??1) z |= 4'b0100; 
	if(x==?20'b111??1???1???0?0??11) z |= 4'b1000; 
	if(x==?20'b?111??1?0????00???11) z |= 4'b0100; 
	if(x==?20'b?1??01?????100??111?) z |= 4'b0100; 
	if(x==?20'b?1???1110?11????1?1?) z |= 4'b0100; 
	if(x==?20'b??????11?111?00???11) z |= 4'b0100; 
	if(x==?20'b?1?1?1?1??11??0??11?) z |= 4'b0100; 
	if(x==?20'b??1?01?????10?0?111?) z |= 4'b0100; 
	if(x==?20'b?11??1101??????01?1?) z |= 4'b1000; 
	if(x==?20'b?1???111???100????11) z |= 4'b0100; 
	if(x==?20'b11???11??1?0?0??1?1?) z |= 4'b1000; 
	if(x==?20'b??1??111???10?0???11) z |= 4'b0100; 
	if(x==?20'b?111??1???1?0?0???11) z |= 4'b0100; 
	if(x==?20'b11???11??1?0??0?1?1?) z |= 4'b1000; 
	if(x==?20'b111??1?????0?00???11) z |= 4'b1000; 
	if(x==?20'b??11?11?0?1??0??1?1?) z |= 4'b0100; 
	if(x==?20'b?????111??1?000??11?) z |= 4'b0100; 
	if(x==?20'b??11?11?0?1???0?1?1?) z |= 4'b0100; 
	if(x==?20'b11???1??111???0???11) z |= 4'b1000; 
	if(x==?20'b111??11?111????????1) z |= 4'b1000; 
	if(x==?20'b?11?????11???000?1?1) z |= 4'b1000; 
	if(x==?20'b11???110?1???0??1?1?) z |= 4'b1000; 
	if(x==?20'b?1110???1????0??11?1) z |= 4'b0100; 
	if(x==?20'b1????10?1?01????11??) z |= 4'b1000; 
	if(x==?20'b?1110?1??????00???11) z |= 4'b0100; 
	if(x==?20'b?11?011????10???1?1?) z |= 4'b0100; 
	if(x==?20'b11???110?1????0?1?1?) z |= 4'b1000; 
	if(x==?20'b???1?01?10?1????11??) z |= 4'b0100; 
	if(x==?20'b111??1?0?????00???11) z |= 4'b1000; 
	if(x==?20'b??1?01??00???1???1?1) z |= 4'b0100; 
	if(x==?20'b??1??1??11???0?11?11) z |= 4'b1000; 
	if(x==?20'b??11??1??111?0????11) z |= 4'b0100; 
	if(x==?20'b???1?111?1???00?1??1) z |= 4'b0100; 
	if(x==?20'b??11011???1??0??1?1?) z |= 4'b0100; 
	if(x==?20'b??11011???1???0?1?1?) z |= 4'b0100; 
	if(x==?20'b?111?11??111???????1) z |= 4'b0100; 
	if(x==?20'b1?1??11??????0001??1) z |= 4'b1000; 
	if(x==?20'b?1?1?11?????000?1??1) z |= 4'b0100; 
	if(x==?20'b?11???11111??0?????1) z |= 4'b0100; 
	if(x==?20'b111????0???1??0?11?1) z |= 4'b1000; 
	if(x==?20'b??1?1?1??1???000?11?) z |= 4'b1000; 
	if(x==?20'b1?1?1?10?????0??111?) z |= 4'b1000; 
	if(x==?20'b?111????????111???11) z |= 4'b0100; 
	if(x==?20'b?11??110?1?0????1?1?) z |= 4'b1000; 
	if(x==?20'b1?????10?100????11??) z |= 4'b1000; 
	if(x==?20'b?11?011?0?1?????1?1?) z |= 4'b0100; 
	if(x==?20'b?11??1?0111???????11) z |= 4'b1000; 
	if(x==?20'b?11???????11000??1?1) z |= 4'b0100; 
	if(x==?20'b??1???1?011??00?1??1) z |= 4'b0100; 
	if(x==?20'b?11?1?1?1??0?0???11?) z |= 4'b1000; 
	if(x==?20'b?1????10??00??1??1?1) z |= 4'b1000; 
	if(x==?20'b??1??1?1?1???000?11?) z |= 4'b1000; 
	if(x==?20'b?1???10??10??0?0?1??) z |= 4'b1000; 
	if(x==?20'b111?111?1?????0???1?) z |= 4'b1000; 
	if(x==?20'b?11?11???111??0????1) z |= 4'b1000; 
	if(x==?20'b?1?101?1??????0?111?) z |= 4'b0100; 
	if(x==?20'b?1???1???110?00?1??1) z |= 4'b1000; 
	if(x==?20'b?11?1????1?0?00?11??) z |= 4'b1000; 
	if(x==?20'b???101??001?????11??) z |= 4'b0100; 
	if(x==?20'b?11?0?11?1?1????1?1?) z |= 4'b0100; 
	if(x==?20'b11????101????0??111?) z |= 4'b1000; 
	if(x==?20'b?1???1?1??1?000??11?) z |= 4'b0100; 
	if(x==?20'b?111??1?????000???11) z |= 4'b0100; 
	if(x==?20'b?11?0?1??111??????11) z |= 4'b0100; 
	if(x==?20'b????111?????111????1) z |= 4'b0010; 
	if(x==?20'b111??????????111??11) z |= 4'b1000; 
	if(x==?20'b1?1?111?1?????0???11) z |= 4'b1000; 
	if(x==?20'b1?1???101?????0?111?) z |= 4'b1000; 
	if(x==?20'b??1??01??01?0?0??1??) z |= 4'b0100; 
	if(x==?20'b11???11??1????001?1?) z |= 4'b1000; 
	if(x==?20'b111??1???????000??11) z |= 4'b1000; 
	if(x==?20'b?11????10?1??00?11??) z |= 4'b0100; 
	if(x==?20'b???1?11???11?00?1??1) z |= 4'b0100; 
	if(x==?20'b??11?11???1?00??1?1?) z |= 4'b0100; 
	if(x==?20'b?11??1?10??1??0??11?) z |= 4'b0100; 
	if(x==?20'b?111?111???1?0????1?) z |= 4'b0100; 
	if(x==?20'b?1??111?111???0???1?) z |= 4'b1000; 
	if(x==?20'b?????111????111???11) z |= 4'b0100; 
	if(x==?20'b??1??111??0??00???11) z |= 4'b1000; 
	if(x==?20'b??1?111?0????00???11) z |= 4'b0100; 
	if(x==?20'b?1??111??0???00???11) z |= 4'b0100; 
	if(x==?20'b?????1?11???000?111?) z |= 4'b0100; 
	if(x==?20'b?1?101?????1?0??111?) z |= 4'b0100; 
	if(x==?20'b?11??11??1?0???01?1?) z |= 4'b1000; 
	if(x==?20'b??1101?????1??0?111?) z |= 4'b0100; 
	if(x==?20'b111??1101???????1?1?) z |= 4'b1000; 
	if(x==?20'b?1?1?111???1?0????11) z |= 4'b0100; 
	if(x==?20'b?11??11?0?1?0???1?1?) z |= 4'b0100; 
	if(x==?20'b????1?1????1?000111?) z |= 4'b1000; 
	if(x==?20'b?????111?????111???1) z |= 4'b0001; 
	if(x==?20'b?1???111???0?00???11) z |= 4'b1000; 
	if(x==?20'b????111??????111??11) z |= 4'b1000; 
	if(x==?20'b????0?1???11?00?1?11) z |= 4'b0100; 
	if(x==?20'b111?1????1???00???11) z |= 4'b1000; 
	if(x==?20'b?11??110?1?????01?1?) z |= 4'b1000; 
	if(x==?20'b??1??111?111?0????1?) z |= 4'b0100; 
	if(x==?20'b11????1?1????0?0111?) z |= 4'b1000; 
	if(x==?20'b?111011????1????1?1?) z |= 4'b0100; 
	if(x==?20'b?11?1?1?1????0?0?11?) z |= 4'b1000; 
	if(x==?20'b1?1???1?1?????00111?) z |= 4'b1000; 
	if(x==?20'b?11???1?11?0?0??1??1) z |= 4'b1000; 
	if(x==?20'b?11?011???1?0???1?1?) z |= 4'b0100; 
	if(x==?20'b?11???1?11?0??0?1??1) z |= 4'b1000; 
	if(x==?20'b1?1?111?11??????1?1?) z |= 4'b1000; 
	if(x==?20'b?????1??11???0001?11) z |= 4'b1000; 
	if(x==?20'b?111???1??1??00???11) z |= 4'b0100; 
	if(x==?20'b111?111??11?????1???) z |= 4'b1000; 
	if(x==?20'b??1??11?11????001??1) z |= 4'b1000; 
	if(x==?20'b?111?111?11?????1???) z |= 4'b0100; 
	if(x==?20'b?1?1?1?????100??111?) z |= 4'b0100; 
	if(x==?20'b??11?1?????10?0?111?) z |= 4'b0100; 
	if(x==?20'b111??11?1??????01?1?) z |= 4'b1000; 
	if(x==?20'b?11??1??0?11?0??1??1) z |= 4'b0100; 
	if(x==?20'b11???10??10??0???1??) z |= 4'b1000; 
	if(x==?20'b?11??1??0?11??0?1??1) z |= 4'b0100; 
	if(x==?20'b?11??1?1???10?0??11?) z |= 4'b0100; 
	if(x==?20'b1?1??10??10???0??1??) z |= 4'b1000; 
	if(x==?20'b??????1???11000?1?11) z |= 4'b0100; 
	if(x==?20'b??1?11??111???0???11) z |= 4'b1000; 
	if(x==?20'b?11???101??????0111?) z |= 4'b1000; 
	if(x==?20'b??1?111??????000??11) z |= 4'b1000; 
	if(x==?20'b?1?1?01??01??0???1??) z |= 4'b0100; 
	if(x==?20'b?111?11????10???1?1?) z |= 4'b0100; 
	if(x==?20'b?1?1?111??11????1?1?) z |= 4'b0100; 
	if(x==?20'b??11?01??01???0??1??) z |= 4'b0100; 
	if(x==?20'b?1???111????000???11) z |= 4'b0100; 
	if(x==?20'b??11???1???1?00?1?11) z |= 4'b0100; 
	if(x==?20'b?1???11?11?0?0??1?1?) z |= 4'b1000; 
	if(x==?20'b?1???11?11?0??0?1?1?) z |= 4'b1000; 
	if(x==?20'b?1??1?1?1?1??1?1?1??) z |= 4'b1000; 
	if(x==?20'b?1????11?111?0????11) z |= 4'b0100; 
	if(x==?20'b????1?1??100?1??11??) z |= 4'b1000; 
	if(x==?20'b?11?01?????10???111?) z |= 4'b0100; 
	if(x==?20'b?1??1?1??1?1?1?1?1??) z |= 4'b1000; 
	if(x==?20'b?1???1?11?1??1?1?1??) z |= 4'b1000; 
	if(x==?20'b?1???11011???0??1?1?) z |= 4'b1000; 
	if(x==?20'b??11??11?1???00?1?1?) z |= 4'b0100; 
	if(x==?20'b111??11??1?0????1?1?) z |= 4'b1000; 
	if(x==?20'b??1?1?1??1?11?1??1??) z |= 4'b0100; 
	if(x==?20'b?1???11011????0?1?1?) z |= 4'b1000; 
	if(x==?20'b??1??1?11?1?1?1??1??) z |= 4'b0100; 
	if(x==?20'b?11?11???10??0??1?1?) z |= 4'b1000; 
	if(x==?20'b?111?11?0?1?????1?1?) z |= 4'b0100; 
	if(x==?20'b11??11????1??00?1?1?) z |= 4'b1000; 
	if(x==?20'b?11?11???10???0?1?1?) z |= 4'b1000; 
	if(x==?20'b??1??11?0?11?0??1?1?) z |= 4'b0100; 
	if(x==?20'b??1??11?0?11??0?1?1?) z |= 4'b0100; 
	if(x==?20'b??1??1?1?1?11?1??1??) z |= 4'b0100; 
	if(x==?20'b?????1?1001??1??11??) z |= 4'b0100; 
	if(x==?20'b111??110?1??????1?1?) z |= 4'b1000; 
	if(x==?20'b??1??11?1????0001??1) z |= 4'b1000; 
	if(x==?20'b????1?1??100??1?11??) z |= 4'b1000; 
	if(x==?20'b??1?1?101????0??111?) z |= 4'b1000; 
	if(x==?20'b?11???11?01??0??1?1?) z |= 4'b0100; 
	if(x==?20'b?111011???1?????1?1?) z |= 4'b0100; 
	if(x==?20'b?11???11?01???0?1?1?) z |= 4'b0100; 
	if(x==?20'b??1?011???11?0??1?1?) z |= 4'b0100; 
	if(x==?20'b??1?011???11??0?1?1?) z |= 4'b0100; 
	if(x==?20'b?11?1?1111??????1??1) z |= 4'b1000; 
	if(x==?20'b?1???11????1000?1??1) z |= 4'b0100; 
	if(x==?20'b?11?1???1?????001?11) z |= 4'b1000; 
	if(x==?20'b?????1?1001???1?11??) z |= 4'b0100; 
	if(x==?20'b?1???11111???00?1?1?) z |= 4'b1100; 
	if(x==?20'b1???11?01??????01??1) z |= 4'b1000; 
	if(x==?20'b???1??11?0?10???1??1) z |= 4'b0100; 
	if(x==?20'b?1???11?11????001?1?) z |= 4'b1000; 
	if(x==?20'b?11??10??10????0?1??) z |= 4'b1000; 
	if(x==?20'b???1??1???11?00?1?11) z |= 4'b0100; 
	if(x==?20'b?1??01?1???1??0?111?) z |= 4'b0100; 
	if(x==?20'b?1110???00????????11) z |= 4'b0100; 
	if(x==?20'b111????0??00??????11) z |= 4'b1000; 
	if(x==?20'b111???101???????111?) z |= 4'b1000; 
	if(x==?20'b111??11??1?????01?1?) z |= 4'b1000; 
	if(x==?20'b?11??01??01?0????1??) z |= 4'b0100; 
	if(x==?20'b1?1?111??????00???11) z |= 4'b1000; 
	if(x==?20'b1?1???10?????00?111?) z |= 4'b1000; 
	if(x==?20'b??1?111???11?00?1?1?) z |= 4'b1100; 
	if(x==?20'b?1?101???????00?111?) z |= 4'b0100; 
	if(x==?20'b???10?11???10???1??1) z |= 4'b0100; 
	if(x==?20'b1?1?11???10????0?1??) z |= 4'b1000; 
	if(x==?20'b?11?11?1??11????1??1) z |= 4'b0100; 
	if(x==?20'b?1?1?111?????00???11) z |= 4'b0100; 
	if(x==?20'b?111?11???1?0???1?1?) z |= 4'b0100; 
	if(x==?20'b??1??11???1100??1?1?) z |= 4'b0100; 
	if(x==?20'b?11?111?111???????1?) z |= 4'b1000; 
	if(x==?20'b??11???1??1??00?1?11) z |= 4'b0100; 
	if(x==?20'b?11??111??0??0????11) z |= 4'b1000; 
	if(x==?20'b?11?111?0????0????11) z |= 4'b0100; 
	if(x==?20'b1????10??10???0??11?) z |= 4'b1000; 
	if(x==?20'b??1???1?1??0?00??111) z |= 4'b1000; 
	if(x==?20'b?11?111??0????0???11) z |= 4'b0100; 
	if(x==?20'b?11???11?1??00??1?1?) z |= 4'b0100; 
	if(x==?20'b1?1?11???1?0???0?1??) z |= 4'b1000; 
	if(x==?20'b?11101?????1????111?) z |= 4'b0100; 
	if(x==?20'b??1?01101?0?????1??1) z |= 4'b1100; 
	if(x==?20'b???1?01??01??0???11?) z |= 4'b0100; 
	if(x==?20'b?1?1??110?1?0????1??) z |= 4'b0100; 
	if(x==?20'b?1?1??11?01?0????1??) z |= 4'b0100; 
	if(x==?20'b11???1??110????0?1??) z |= 4'b1000; 
	if(x==?20'b?1??1?1??11??1?1?1??) z |= 4'b1000; 
	if(x==?20'b?11?11????1???001?1?) z |= 4'b1000; 
	if(x==?20'b????1?1?1?1?1?1??1??) z |= 4'b0010; 
	if(x==?20'b?11??111???0??0???11) z |= 4'b1000; 
	if(x==?20'b??1?1?1??11?1?1??1??) z |= 4'b0100; 
	if(x==?20'b????11??11??11??1???) z |= 4'b0010; 
	if(x==?20'b?1???1??0??1?00??111) z |= 4'b0100; 
	if(x==?20'b?1???1?1?11??1?1?1??) z |= 4'b1000; 
	if(x==?20'b?11??111?111??????1?) z |= 4'b0100; 
	if(x==?20'b?11?1???11???00?1??1) z |= 4'b1000; 
	if(x==?20'b??1??1?1?11?1?1??1??) z |= 4'b0100; 
	if(x==?20'b1?1??11?1????00?1??1) z |= 4'b1000; 
	if(x==?20'b?11?1?1??????000?11?) z |= 4'b1000; 
	if(x==?20'b?????1?1?1?1?1?1?1??) z |= 4'b0001; 
	if(x==?20'b??1??1??11????001?11) z |= 4'b1000; 
	if(x==?20'b?1???11?01???00??11?) z |= 4'b0100; 
	if(x==?20'b?11??1?1????000??11?) z |= 4'b0100; 
	if(x==?20'b?1???10?110??0???1??) z |= 4'b1000; 
	if(x==?20'b??1??11??1???0001??1) z |= 4'b1000; 
	if(x==?20'b??11??1??0110????1??) z |= 4'b0100; 
	if(x==?20'b?1?1?11????1?00?1??1) z |= 4'b0100; 
	if(x==?20'b???1??110??10???11??) z |= 4'b0100; 
	if(x==?20'b??1??11???10?00??11?) z |= 4'b1000; 
	if(x==?20'b?1???11???1?000?1??1) z |= 4'b0100; 
	if(x==?20'b11???11?11???0??1?1?) z |= 4'b1000; 
	if(x==?20'b11???11?11????0?1?1?) z |= 4'b1000; 
	if(x==?20'b111??1??1????00???11) z |= 4'b1000; 
	if(x==?20'b111??10??10??????1??) z |= 4'b1000; 
	if(x==?20'b?11????1??11?00?1??1) z |= 4'b0100; 
	if(x==?20'b?11?1????1????001?11) z |= 4'b1000; 
	if(x==?20'b?11?111??????0?0??11) z |= 4'b1000; 
	if(x==?20'b???1??1?0101?????11?) z |= 4'b0100; 
	if(x==?20'b1???11?0?1?????01??1) z |= 4'b1000; 
	if(x==?20'b?11?11???????0001?1?) z |= 4'b1000; 
	if(x==?20'b?111?01??01??????1??) z |= 4'b0100; 
	if(x==?20'b?111??1????1?00???11) z |= 4'b0100; 
	if(x==?20'b?11???11????000?1?1?) z |= 4'b0100; 
	if(x==?20'b?11??111????0?0???11) z |= 4'b0100; 
	if(x==?20'b??????1110??10??11??) z |= 4'b0100; 
	if(x==?20'b1???1?10?10?????11??) z |= 4'b1000; 
	if(x==?20'b??1??01??011??0??1??) z |= 4'b0100; 
	if(x==?20'b1????1??1010?????11?) z |= 4'b1000; 
	if(x==?20'b1?1?1??0?1?????0?1?1) z |= 4'b1000; 
	if(x==?20'b???10?11??1?0???1??1) z |= 4'b0100; 
	if(x==?20'b?1???1??111??00???11) z |= 4'b1000; 
	if(x==?20'b??11?11???11?0??1?1?) z |= 4'b0100; 
	if(x==?20'b??11?11???11??0?1?1?) z |= 4'b0100; 
	if(x==?20'b?11?0??1?????00?1?11) z |= 4'b0100; 
	if(x==?20'b?11?0???1????00?11?1) z |= 4'b0100; 
	if(x==?20'b1???1?10?????0?0?1?1) z |= 4'b1000; 
	if(x==?20'b?1?10??1??1?0????1?1) z |= 4'b0100; 
	if(x==?20'b??1???1??111?00???11) z |= 4'b0100; 
	if(x==?20'b??????11??11??111???) z |= 4'b0001; 
	if(x==?20'b11?????011?????0?1?1) z |= 4'b1000; 
	if(x==?20'b???101?1?01?????11??) z |= 4'b0100; 
	if(x==?20'b??1???11??11?00?1?1?) z |= 4'b0100; 
	if(x==?20'b???101?1????0?0??1?1) z |= 4'b0100; 
	if(x==?20'b????11????01??0111??) z |= 4'b1000; 
	if(x==?20'b??110???00??????1?11) z |= 4'b0100; 
	if(x==?20'b?1???11???1?000??11?) z |= 4'b0100; 
	if(x==?20'b11?????0??00????1?11) z |= 4'b1000; 
	if(x==?20'b?11????0???1?00?11?1) z |= 4'b1000; 
	if(x==?20'b1?1???1??1???1?1?1?1) z |= 4'b1000; 
	if(x==?20'b1????1??110????0?11?) z |= 4'b1000; 
	if(x==?20'b????11???11?11??1???) z |= 4'b0010; 
	if(x==?20'b1?1??11??1???00?1??1) z |= 4'b1000; 
	if(x==?20'b??110?????110????1?1) z |= 4'b0100; 
	if(x==?20'b???1??11??1?01???11?) z |= 4'b0100; 
	if(x==?20'b?11?1????????0001?11) z |= 4'b1000; 
	if(x==?20'b?1?1?1????1?1?1??1?1) z |= 4'b0100; 
	if(x==?20'b?11??11?11?????01?1?) z |= 4'b1000; 
	if(x==?20'b??1?111?1????00???11) z |= 4'b1000; 
	if(x==?20'b??1???101????00?111?) z |= 4'b1000; 
	if(x==?20'b?11????1????000?1?11) z |= 4'b0100; 
	if(x==?20'b?11?????1???000?11?1) z |= 4'b0100; 
	if(x==?20'b?1?1?11???1??00?1??1) z |= 4'b0100; 
	if(x==?20'b??????11?11?11??1?1?) z |= 4'b0100; 
	if(x==?20'b1???11???1????10?11?) z |= 4'b1000; 
	if(x==?20'b?1?10?1??01??0???1??) z |= 4'b0100; 
	if(x==?20'b??1??01?0???0?0??11?) z |= 4'b0100; 
	if(x==?20'b?11????????1?00011?1) z |= 4'b1000; 
	if(x==?20'b?1??01?????1?00?111?) z |= 4'b0100; 
	if(x==?20'b?1???10????0?0?0?11?) z |= 4'b1000; 
	if(x==?20'b???1??1???1101???11?) z |= 4'b0100; 
	if(x==?20'b11???10?1??????011??) z |= 4'b1000; 
	if(x==?20'b?1???111???1?00???11) z |= 4'b0100; 
	if(x==?20'b?11??11???110???1?1?) z |= 4'b0100; 
	if(x==?20'b?1??11??1?10???0?1??) z |= 4'b1000; 
	if(x==?20'b??1????1??11?00?1?11) z |= 4'b0100; 
	if(x==?20'b??1???1101?10????1??) z |= 4'b0100; 
	if(x==?20'b??11?01????10???11??) z |= 4'b0100; 
	if(x==?20'b?1???110?1?0???0?1??) z |= 4'b1000; 
	if(x==?20'b??1?011?0?1?0????1??) z |= 4'b0100; 
	if(x==?20'b??????11?11???111???) z |= 4'b0001; 
	if(x==?20'b????11???11???111?1?) z |= 4'b1000; 
	if(x==?20'b?1??111??1???1?1?1??) z |= 4'b1000; 
	if(x==?20'b?1?1?01?01??????11??) z |= 4'b0100; 
	if(x==?20'b111?1????????00?1?11) z |= 4'b1000; 
	if(x==?20'b?1?1??1??1??1?1??11?) z |= 4'b0100; 
	if(x==?20'b?1???11?1?1??1?1?1??) z |= 4'b1000; 
	if(x==?20'b????11?011?????01??1) z |= 4'b1000; 
	if(x==?20'b111??11?11??????1?1?) z |= 4'b1000; 
	if(x==?20'b11???11??1???00?1?1?) z |= 4'b1000; 
	if(x==?20'b???1011??0?1????1??1) z |= 4'b0100; 
	if(x==?20'b1?1??1????1??1?1?11?) z |= 4'b1000; 
	if(x==?20'b11??11??110??????1??) z |= 4'b1000; 
	if(x==?20'b??1??11??1?11?1??1??) z |= 4'b0100; 
	if(x==?20'b?1?1?01?0????0???11?) z |= 4'b0100; 
	if(x==?20'b??11?11???1??00?1?1?) z |= 4'b0100; 
	if(x==?20'b1???111??????1?01??1) z |= 4'b1000; 
	if(x==?20'b111?1?????00??????11) z |= 4'b1000; 
	if(x==?20'b?11??11??1?0?0??1?1?) z |= 4'b1000; 
	if(x==?20'b1????1?0?10???0??11?) z |= 4'b1000; 
	if(x==?20'b??11?11?01???1???1??) z |= 4'b0100; 
	if(x==?20'b?11??11??1?0??0?1?1?) z |= 4'b1000; 
	if(x==?20'b????1?101????0?0?1?1) z |= 4'b1000; 
	if(x==?20'b1?1??10????0??0??11?) z |= 4'b1000; 
	if(x==?20'b?11??11?0?1??0??1?1?) z |= 4'b0100; 
	if(x==?20'b?111???100????????11) z |= 4'b0100; 
	if(x==?20'b?11??11?0?1???0?1?1?) z |= 4'b0100; 
	if(x==?20'b?11??1??111???0???11) z |= 4'b1000; 
	if(x==?20'b?111?11???11????1?1?) z |= 4'b0100; 
	if(x==?20'b????0?11??110???1??1) z |= 4'b0100; 
	if(x==?20'b?1?11?1?1?1??1???1??) z |= 4'b0100; 
	if(x==?20'b???10?1??01??0???11?) z |= 4'b0100; 
	if(x==?20'b111?1??0??0???????11) z |= 4'b1000; 
	if(x==?20'b111?????1?00??????11) z |= 4'b1000; 
	if(x==?20'b?1?11?1??1?1?1???1??) z |= 4'b0100; 
	if(x==?20'b?1?1?1?11?1??1???1??) z |= 4'b0100; 
	if(x==?20'b?11???1??111?0????11) z |= 4'b0100; 
	if(x==?20'b1?1???1?1????00?111?) z |= 4'b1000; 
	if(x==?20'b?1??1?10?10???0??1??) z |= 4'b1000; 
	if(x==?20'b????11??11???11?1???) z |= 4'b0010; 
	if(x==?20'b??11??11?011?????1??) z |= 4'b0100; 
	if(x==?20'b1???11??1??1???01??1) z |= 4'b1000; 
	if(x==?20'b?1110??1?0????????11) z |= 4'b0100; 
	if(x==?20'b?1?1?1?1?1?1?1???1??) z |= 4'b0100; 
	if(x==?20'b???1?111????0?1?1??1) z |= 4'b0100; 
	if(x==?20'b??????11?0??0?1?1?11) z |= 4'b0100; 
	if(x==?20'b????01?1???10?0??1?1) z |= 4'b0100; 
	if(x==?20'b1?1?1?1?1?1???1??1??) z |= 4'b1000; 
	if(x==?20'b?111????00?1??????11) z |= 4'b0100; 
	if(x==?20'b??1???10?100????11??) z |= 4'b1000; 
	if(x==?20'b?1?1??11?0??0???1??1) z |= 4'b0100; 
	if(x==?20'b1?1?1?1??1?1??1??1??) z |= 4'b1000; 
	if(x==?20'b111??11?1????0??1?1?) z |= 4'b1000; 
	if(x==?20'b11???11???10??1??1??) z |= 4'b1000; 
	if(x==?20'b1?1??1?11?1???1??1??) z |= 4'b1000; 
	if(x==?20'b?1?1?1?????1?00?111?) z |= 4'b0100; 
	if(x==?20'b??1?01?1?01??0???1??) z |= 4'b0100; 
	if(x==?20'b111??11?1?????0?1?1?) z |= 4'b1000; 
	if(x==?20'b???????11001????111?) z |= 4'b0100; 
	if(x==?20'b????11??11????10?11?) z |= 4'b1000; 
	if(x==?20'b1?1??1?1?1?1??1??1??) z |= 4'b1000; 
	if(x==?20'b?1??01??001?????11??) z |= 4'b0100; 
	if(x==?20'b??????11??11?11?1???) z |= 4'b0001; 
	if(x==?20'b??????11??1101???11?) z |= 4'b0100; 
	if(x==?20'b????0?11????0?1?1?11) z |= 4'b0100; 
	if(x==?20'b?11???101????0??111?) z |= 4'b1000; 
	if(x==?20'b1?1?11?0???????01??1) z |= 4'b1000; 
	if(x==?20'b?11??11??1????001?1?) z |= 4'b1000; 
	if(x==?20'b1???11?011??????1??1) z |= 4'b1000; 
	if(x==?20'b?1?10?11????0???1??1) z |= 4'b0100; 
	if(x==?20'b????11????01?10?11??) z |= 4'b1000; 
	if(x==?20'b?111?11????1?0??1?1?) z |= 4'b0100; 
	if(x==?20'b?1???11???11?00?1??1) z |= 4'b0100; 
	if(x==?20'b11??11??1?1????0?1??) z |= 4'b1000; 
	if(x==?20'b?111?11????1??0?1?1?) z |= 4'b0100; 
	if(x==?20'b?11??11???1?00??1?1?) z |= 4'b0100; 
	if(x==?20'b????1??011?0????1?11) z |= 4'b1000; 
	if(x==?20'b1?1?1??011???????1?1) z |= 4'b1000; 
	if(x==?20'b?1???11??11??1?1?1??) z |= 4'b1000; 
	if(x==?20'b????1???1001????111?) z |= 4'b1010; 
	if(x==?20'b?????11?11??11??1???) z |= 4'b0010; 
	if(x==?20'b??1??11??11?1?1??1??) z |= 4'b0100; 
	if(x==?20'b??11??11?1?10????1??) z |= 4'b0100; 
	if(x==?20'b??????1110???01?11??) z |= 4'b0100; 
	if(x==?20'b?11??11?1?1??00?1?1?) z |= 4'b1100; 
	if(x==?20'b?11?01?????1??0?111?) z |= 4'b0100; 
	if(x==?20'b?11??11??1?1?00?1?1?) z |= 4'b1100; 
	if(x==?20'b1???111??1????00???1) z |= 4'b1000; 
	if(x==?20'b???10?11??11????1??1) z |= 4'b0100; 
	if(x==?20'b1?1?1???0??0?????111) z |= 4'b1000; 
	if(x==?20'b?1?1??110???0????11?) z |= 4'b0100; 
	if(x==?20'b1?1?111?1??0???????1) z |= 4'b1000; 
	if(x==?20'b?11???1?1????0?0111?) z |= 4'b1000; 
	if(x==?20'b????0??10?11????1?11) z |= 4'b0100; 
	if(x==?20'b111??1???10????0?1??) z |= 4'b1000; 
	if(x==?20'b1?1?11?????0???0?11?) z |= 4'b1000; 
	if(x==?20'b??11??11011??????1??) z |= 4'b0100; 
	if(x==?20'b?1?1???10??0?????111) z |= 4'b0100; 
	if(x==?20'b???1?111??1?00?????1) z |= 4'b0100; 
	if(x==?20'b11??11???110?????1??) z |= 4'b1000; 
	if(x==?20'b?1?11?1??11??1???1??) z |= 4'b0100; 
	if(x==?20'b?1?10??1??11?????1?1) z |= 4'b0100; 
	if(x==?20'b1???1?1?110?????11??) z |= 4'b1000; 
	if(x==?20'b?111??1??01?0????1??) z |= 4'b0100; 
	if(x==?20'b1?1?1???11?????0?1?1) z |= 4'b1000; 
	if(x==?20'b?1?1?1110??1???????1) z |= 4'b0100; 
	if(x==?20'b?1?1?1?1?11??1???1??) z |= 4'b0100; 
	if(x==?20'b1?1??1??1??0???0?11?) z |= 4'b1000; 
	if(x==?20'b?11??1?????10?0?111?) z |= 4'b0100; 
	if(x==?20'b????11111111??????1?) z |= 4'b1100; 
	if(x==?20'b11??1?????00????1?11) z |= 4'b1000; 
	if(x==?20'b1???11?01????0??1??1) z |= 4'b1000; 
	if(x==?20'b1??????0?1???0?0?111) z |= 4'b1000; 
	if(x==?20'b???1??11?0?1?0??1??1) z |= 4'b0100; 
	if(x==?20'b?1?1??1?0??10????11?) z |= 4'b0100; 
	if(x==?20'b1???11?01?????0?1??1) z |= 4'b1000; 
	if(x==?20'b?11??10??10??0???1??) z |= 4'b1000; 
	if(x==?20'b????11???11??11?1???) z |= 4'b0010; 
	if(x==?20'b1???1?1?1????0?0?1?1) z |= 4'b1000; 
	if(x==?20'b???1??11?0?1??0?1??1) z |= 4'b0100; 
	if(x==?20'b1?1?1?1??11???1??1??) z |= 4'b1000; 
	if(x==?20'b??11???100??????1?11) z |= 4'b0100; 
	if(x==?20'b??????11?11??11?1???) z |= 4'b0001; 
	if(x==?20'b????11???11??11?1?1?) z |= 4'b1000; 
	if(x==?20'b???10?????1?0?0??111) z |= 4'b0100; 
	if(x==?20'b?1???10?1?0???0??11?) z |= 4'b1000; 
	if(x==?20'b111??11??1???0??1?1?) z |= 4'b1000; 
	if(x==?20'b1?1??1?1?11???1??1??) z |= 4'b1000; 
	if(x==?20'b??????11?11??11?1?1?) z |= 4'b0100; 
	if(x==?20'b????11?0?1????001??1) z |= 4'b1000; 
	if(x==?20'b111??11??1????0?1?1?) z |= 4'b1000; 
	if(x==?20'b?11??01??01???0??1??) z |= 4'b0100; 
	if(x==?20'b11??????1?00????1?11) z |= 4'b1000; 
	if(x==?20'b1????110?1?0????11??) z |= 4'b1000; 
	if(x==?20'b11??1?1??10???0??1??) z |= 4'b1000; 
	if(x==?20'b1?1?11???10??0???1??) z |= 4'b1000; 
	if(x==?20'b???10?11???1?0??1??1) z |= 4'b0100; 
	if(x==?20'b???1011?0?1?????11??) z |= 4'b0100; 
	if(x==?20'b?1?1???1??110????1?1) z |= 4'b0100; 
	if(x==?20'b???10?11???1??0?1??1) z |= 4'b0100; 
	if(x==?20'b?111?11???1??0??1?1?) z |= 4'b0100; 
	if(x==?20'b?????11???11??111???) z |= 4'b0001; 
	if(x==?20'b????0?11??1?00??1??1) z |= 4'b0100; 
	if(x==?20'b??110??1?0??????1?11) z |= 4'b0100; 
	if(x==?20'b?111?11???1???0?1?1?) z |= 4'b0100; 
	if(x==?20'b???1?1?1?011????11??) z |= 4'b0100; 
	if(x==?20'b??1??01??0?1?0???11?) z |= 4'b0100; 
	if(x==?20'b1?1?11???1?0?0???1??) z |= 4'b1000; 
	if(x==?20'b???1?1?1???10?0??1?1) z |= 4'b0100; 
	if(x==?20'b?1???10?1?0???0?11??) z |= 4'b1000; 
	if(x==?20'b??11????00?1????1?11) z |= 4'b0100; 
	if(x==?20'b1?1?11???1?0??0??1??) z |= 4'b1000; 
	if(x==?20'b?11???11?1???00?1?1?) z |= 4'b0100; 
	if(x==?20'b11????1??100????11??) z |= 4'b1000; 
	if(x==?20'b11???1??110??0???1??) z |= 4'b1000; 
	if(x==?20'b?1?1??110?1??0???1??) z |= 4'b0100; 
	if(x==?20'b?11?11????1??00?1?1?) z |= 4'b1000; 
	if(x==?20'b?1?1??110?1???0??1??) z |= 4'b0100; 
	if(x==?20'b?1?1??11?01???0??1??) z |= 4'b0100; 
	if(x==?20'b1???11??1?????001??1) z |= 4'b1000; 
	if(x==?20'b??11?1?1?01??0???1??) z |= 4'b0100; 
	if(x==?20'b??1??1110???00?????1) z |= 4'b0100; 
	if(x==?20'b?1???1101?10?????1??) z |= 4'b1000; 
	if(x==?20'b1???11??1?0??0??11??) z |= 4'b1000; 
	if(x==?20'b??1?011?01?1?????1??) z |= 4'b0100; 
	if(x==?20'b?1??111????0??00???1) z |= 4'b1000; 
	if(x==?20'b??11?1??001?????11??) z |= 4'b0100; 
	if(x==?20'b1?1?1?1????1???111??) z |= 4'b1000; 
	if(x==?20'b??1??01??0?1?0??11??) z |= 4'b0100; 
	if(x==?20'b1????110?1?????0?11?) z |= 4'b1000; 
	if(x==?20'b???1??11????0?1?1?11) z |= 4'b0100; 
	if(x==?20'b?????11??11?11??1???) z |= 4'b0010; 
	if(x==?20'b11???1??11?0??0??1??) z |= 4'b1000; 
	if(x==?20'b???1?01?????0?0?111?) z |= 4'b0100; 
	if(x==?20'b?1??1????100??0?11??) z |= 4'b1000; 
	if(x==?20'b1????10??????0?0111?) z |= 4'b1000; 
	if(x==?20'b?1?10?1?01??????11??) z |= 4'b0100; 
	if(x==?20'b???1011???1?0????11?) z |= 4'b0100; 
	if(x==?20'b???1??11???100??1??1) z |= 4'b0100; 
	if(x==?20'b?????111???10?1?1??1) z |= 4'b0100; 
	if(x==?20'b1???1???11?0????1?11) z |= 4'b1000; 
	if(x==?20'b??1????1001??0??11??) z |= 4'b0100; 
	if(x==?20'b??11??1??011?0???1??) z |= 4'b0100; 
	if(x==?20'b1???111?1??0??????11) z |= 4'b1000; 
	if(x==?20'b??11??1??011??0??1??) z |= 4'b0100; 
	if(x==?20'b??1?11?01??????01??1) z |= 4'b1000; 
	if(x==?20'b?1???10?1????0?0?11?) z |= 4'b1000; 
	if(x==?20'b?1????11?0?10???1??1) z |= 4'b0100; 
	if(x==?20'b????111?00???0????11) z |= 4'b0100; 
	if(x==?20'b?1???110?????1?01??1) z |= 4'b1000; 
	if(x==?20'b?1????1???11?00?1?11) z |= 4'b0100; 
	if(x==?20'b?????111??00??0???11) z |= 4'b1000; 
	if(x==?20'b???1?1110??1??????11) z |= 4'b0100; 
	if(x==?20'b??1??01????10?0??11?) z |= 4'b0100; 
	if(x==?20'b1???11?0?1???0??1??1) z |= 4'b1000; 
	if(x==?20'b1???11?0?1????0?1??1) z |= 4'b1000; 
	if(x==?20'b???1???10?11????1?11) z |= 4'b0100; 
	if(x==?20'b????11?0?????0?11?11) z |= 4'b1000; 
	if(x==?20'b?1?1??1???1?01???11?) z |= 4'b0100; 
	if(x==?20'b?1??0?11???10???1??1) z |= 4'b0100; 
	if(x==?20'b?1?10?1?0????0???11?) z |= 4'b0100; 
	if(x==?20'b?????11??11???111???) z |= 4'b0001; 
	if(x==?20'b1?1?1??0?1???0???1?1) z |= 4'b1000; 
	if(x==?20'b???10?11??1??0??1??1) z |= 4'b0100; 
	if(x==?20'b????111?11????00???1) z |= 4'b1000; 
	if(x==?20'b???10?11??1???0?1??1) z |= 4'b0100; 
	if(x==?20'b??1?011?????0?1?1??1) z |= 4'b0100; 
	if(x==?20'b?1??1????10???0011??) z |= 4'b1000; 
	if(x==?20'b?11???11?100????11??) z |= 4'b1100; 
	if(x==?20'b1?1??1?0???0??0??11?) z |= 4'b1000; 
	if(x==?20'b?1???01??01??0???11?) z |= 4'b0100; 
	if(x==?20'b1?1??1???1????10?11?) z |= 4'b1000; 
	if(x==?20'b?11??1??110????0?1??) z |= 4'b1000; 
	if(x==?20'b?1??11??1110?????1??) z |= 4'b1000; 
	if(x==?20'b11?????011???0???1?1) z |= 4'b1000; 
	if(x==?20'b?1?10??1??1???0??1?1) z |= 4'b0100; 
	if(x==?20'b11?????011????0??1?1) z |= 4'b1000; 
	if(x==?20'b?11?0??01??1?????111) z |= 4'b1100; 
	if(x==?20'b??1?011?0???0????11?) z |= 4'b0100; 
	if(x==?20'b??1????1?01?00??11??) z |= 4'b0100; 
	if(x==?20'b????111???0??0?0??11) z |= 4'b1000; 
	if(x==?20'b??1???110111?????1??) z |= 4'b0100; 
	if(x==?20'b1???11???1????001??1) z |= 4'b1000; 
	if(x==?20'b?11??11??11??11?1???) z |= 4'b1100; 
	if(x==?20'b?1???110???0???0?11?) z |= 4'b1000; 
	if(x==?20'b?????111??1100?????1) z |= 4'b0100; 
	if(x==?20'b1????1??110???0??11?) z |= 4'b1000; 
	if(x==?20'b???????011???0?0?111) z |= 4'b1000; 
	if(x==?20'b1?1?1????1???0?0?1?1) z |= 4'b1000; 
	if(x==?20'b1????1101??1????1??1) z |= 4'b1000; 
	if(x==?20'b??11??1?011??0???1??) z |= 4'b0100; 
	if(x==?20'b1???1?10?1????0??11?) z |= 4'b1000; 
	if(x==?20'b???1??11??1?00??1??1) z |= 4'b0100; 
	if(x==?20'b?11???1??0110????1??) z |= 4'b0100; 
	if(x==?20'b?????1110???00????11) z |= 4'b0100; 
	if(x==?20'b??110?????11?0???1?1) z |= 4'b0100; 
	if(x==?20'b????111????0??00??11) z |= 4'b1000; 
	if(x==?20'b?????111?0??0?0???11) z |= 4'b0100; 
	if(x==?20'b?????111??1?0?1?1??1) z |= 4'b0100; 
	if(x==?20'b??110?????11??0??1?1) z |= 4'b0100; 
	if(x==?20'b???1??11??1??10??11?) z |= 4'b0100; 
	if(x==?20'b?1????110??10???11??) z |= 4'b0100; 
	if(x==?20'b111?1???1?0???????11) z |= 4'b1000; 
	if(x==?20'b1?1?1110?1???????1??) z |= 4'b1000; 
	if(x==?20'b?11??11?11???0??1?1?) z |= 4'b1000; 
	if(x==?20'b1?1?11?01???????1??1) z |= 4'b1000; 
	if(x==?20'b11???1???110??0??1??) z |= 4'b1000; 
	if(x==?20'b?11??11?11????0?1?1?) z |= 4'b1000; 
	if(x==?20'b?1?1??11?0?1????1??1) z |= 4'b0100; 
	if(x==?20'b1???11???1???01??11?) z |= 4'b1000; 
	if(x==?20'b?1?1?111??1??1???1??) z |= 4'b0100; 
	if(x==?20'b?1??1?1?110???0??1??) z |= 4'b1000; 
	if(x==?20'b?1?1???1??1?0?0??1?1) z |= 4'b0100; 
	if(x==?20'b???101?1??1??0???11?) z |= 4'b0100; 
	if(x==?20'b1?1?111??1????1??1??) z |= 4'b1000; 
	if(x==?20'b??1?11?0?1?????01??1) z |= 4'b1000; 
	if(x==?20'b?1????1?0101?????11?) z |= 4'b0100; 
	if(x==?20'b1???111?1??0????11??) z |= 4'b1000; 
	if(x==?20'b???1??1??011?0???11?) z |= 4'b0100; 
	if(x==?20'b11??1?????????10111?) z |= 4'b1000; 
	if(x==?20'b????0?????110?0??111) z |= 4'b0100; 
	if(x==?20'b?1?10111??1??????1??) z |= 4'b0100; 
	if(x==?20'b?1?1?11?1?1??1???1??) z |= 4'b0100; 
	if(x==?20'b11???11011???????1??) z |= 4'b1000; 
	if(x==?20'b??1?1?10?10?????11??) z |= 4'b1000; 
	if(x==?20'b??1??1??1010?????11?) z |= 4'b1000; 
	if(x==?20'b??11???1????0?1?111?) z |= 4'b0100; 
	if(x==?20'b?1?10?11???1????1??1) z |= 4'b0100; 
	if(x==?20'b11???10?1????0??11??) z |= 4'b1000; 
	if(x==?20'b?1110?1?0?????????11) z |= 4'b0100; 
	if(x==?20'b1????1??11???01??11?) z |= 4'b1000; 
	if(x==?20'b?1????1?1100????11??) z |= 4'b1000; 
	if(x==?20'b?1?1?11??1?1?1???1??) z |= 4'b0100; 
	if(x==?20'b?1??0?11??1?0???1??1) z |= 4'b0100; 
	if(x==?20'b???1??1???11?10??11?) z |= 4'b0100; 
	if(x==?20'b?????11?11???11?1???) z |= 4'b0010; 
	if(x==?20'b11???1101?1??????1??) z |= 4'b1000; 
	if(x==?20'b?11??11???11?0??1?1?) z |= 4'b0100; 
	if(x==?20'b?1??11??1?10?0???1??) z |= 4'b1000; 
	if(x==?20'b?111???1?0?1??????11) z |= 4'b0100; 
	if(x==?20'b11??111???????00???1) z |= 4'b1000; 
	if(x==?20'b?11??11???11??0?1?1?) z |= 4'b0100; 
	if(x==?20'b1???111?11????0????1) z |= 4'b1000; 
	if(x==?20'b1???11???1???0?0?11?) z |= 4'b1000; 
	if(x==?20'b???1?111?0?1????11??) z |= 4'b0100; 
	if(x==?20'b??11?111????00?????1) z |= 4'b0100; 
	if(x==?20'b111??1?0???0??????11) z |= 4'b1000; 
	if(x==?20'b??1?01?101??????11??) z |= 4'b0100; 
	if(x==?20'b??11011??1?1?????1??) z |= 4'b0100; 
	if(x==?20'b??1???1101?1??0??1??) z |= 4'b0100; 
	if(x==?20'b?????11011?????0?11?) z |= 4'b1000; 
	if(x==?20'b??1?1?10?????0?0?1?1) z |= 4'b1000; 
	if(x==?20'b?1???110?1?0?0???1??) z |= 4'b1000; 
	if(x==?20'b??11?01????1??0?11??) z |= 4'b0100; 
	if(x==?20'b111??1??110??????1??) z |= 4'b1000; 
	if(x==?20'b1?1?11??1??0?????11?) z |= 4'b1000; 
	if(x==?20'b1?1?11??1??????01??1) z |= 4'b1000; 
	if(x==?20'b?1??1?10??10????11??) z |= 4'b1000; 
	if(x==?20'b1???1???1?0???0?111?) z |= 4'b1000; 
	if(x==?20'b1?1??11?1?1???1??1??) z |= 4'b1000; 
	if(x==?20'b?????10?1????0?0111?) z |= 4'b1000; 
	if(x==?20'b1???11???????0001??1) z |= 4'b1000; 
	if(x==?20'b?11????011?????0?1?1) z |= 4'b1000; 
	if(x==?20'b??1?011?0?1???0??1??) z |= 4'b0100; 
	if(x==?20'b?1?????0?1???000?1?1) z |= 4'b1000; 
	if(x==?20'b?1??01?1?01?????11??) z |= 4'b0100; 
	if(x==?20'b??11011???11?????1??) z |= 4'b0100; 
	if(x==?20'b?1?1????0???0?0??111) z |= 4'b0100; 
	if(x==?20'b???1??11????000?1??1) z |= 4'b0100; 
	if(x==?20'b??1??1?1?011?0???1??) z |= 4'b0100; 
	if(x==?20'b???1??11??1?0?0??11?) z |= 4'b0100; 
	if(x==?20'b1?1????????0?0?0?111) z |= 4'b1000; 
	if(x==?20'b?1??01?1????0?0??1?1) z |= 4'b0100; 
	if(x==?20'b11???11??????1?01??1) z |= 4'b1000; 
	if(x==?20'b?11?0???00??????1?11) z |= 4'b0100; 
	if(x==?20'b?11????0??00????1?11) z |= 4'b1000; 
	if(x==?20'b?????11???11?11?1???) z |= 4'b0001; 
	if(x==?20'b??1?0?????1?000??1?1) z |= 4'b0100; 
	if(x==?20'b??11011?0????????11?) z |= 4'b0100; 
	if(x==?20'b??1??1??0011????11??) z |= 4'b0100; 
	if(x==?20'b?1?1??110??1?????11?) z |= 4'b0100; 
	if(x==?20'b??????11???10?1?1?11) z |= 4'b0100; 
	if(x==?20'b?????01????10?0?111?) z |= 4'b0100; 
	if(x==?20'b1?1?11?????1???01??1) z |= 4'b1000; 
	if(x==?20'b1???11???????0?11?11) z |= 4'b1000; 
	if(x==?20'b??1??1??110????0?11?) z |= 4'b1000; 
	if(x==?20'b11???110???0?????11?) z |= 4'b1000; 
	if(x==?20'b?1?1??11???10???1??1) z |= 4'b0100; 
	if(x==?20'b???1?111??11?0?????1) z |= 4'b0100; 
	if(x==?20'b11?????0?????0?0?111) z |= 4'b1000; 
	if(x==?20'b????011???110????11?) z |= 4'b0100; 
	if(x==?20'b?1??1?10?1?????0?11?) z |= 4'b1000; 
	if(x==?20'b??110???????0?0??111) z |= 4'b0100; 
	if(x==?20'b?11?0?????110????1?1) z |= 4'b0100; 
	if(x==?20'b???1???1?0?1?0??111?) z |= 4'b0100; 
	if(x==?20'b?1????11??1?01???11?) z |= 4'b0100; 
	if(x==?20'b?111??1??011?????1??) z |= 4'b0100; 
	if(x==?20'b???1?1110????0????11) z |= 4'b0100; 
	if(x==?20'b??1?1?1011???0???11?) z |= 4'b1100; 
	if(x==?20'b?1?1?1?11????1??11??) z |= 4'b0100; 
	if(x==?20'b1???111????0??0???11) z |= 4'b1000; 
	if(x==?20'b?1??1?10???0??0??11?) z |= 4'b1000; 
	if(x==?20'b??1?01?10????0???11?) z |= 4'b0100; 
	if(x==?20'b??11?11?????0?1?1??1) z |= 4'b0100; 
	if(x==?20'b????11?011???0??1??1) z |= 4'b1000; 
	if(x==?20'b????11?011????0?1??1) z |= 4'b1000; 
	if(x==?20'b??1?111?00????????11) z |= 4'b0100; 
	if(x==?20'b??1?11???1????10?11?) z |= 4'b1000; 
	if(x==?20'b??1?01?1??1?0????11?) z |= 4'b0100; 
	if(x==?20'b?1???1?01?0???0??11?) z |= 4'b1000; 
	if(x==?20'b?1???111??00??????11) z |= 4'b1000; 
	if(x==?20'b111?11???1?????0?1??) z |= 4'b1000; 
	if(x==?20'b1?1?11?0?1??????1??1) z |= 4'b1000; 
	if(x==?20'b1?1?11??1??????0?11?) z |= 4'b1000; 
	if(x==?20'b11???1??11?0????1??1) z |= 4'b1000; 
	if(x==?20'b?1?1?1?11?????1?11??) z |= 4'b0100; 
	if(x==?20'b?11??10?1??????011??) z |= 4'b1000; 
	if(x==?20'b?1????1???1101???11?) z |= 4'b0100; 
	if(x==?20'b?111??11??1?0????1??) z |= 4'b0100; 
	if(x==?20'b??1?0?1??0?1?0???11?) z |= 4'b0100; 
	if(x==?20'b1?1?1?1????1??1?11??) z |= 4'b1000; 
	if(x==?20'b111?????1111???????1) z |= 4'b1000; 
	if(x==?20'b?1?10?11??1?????1??1) z |= 4'b0100; 
	if(x==?20'b?111????1111???????1) z |= 4'b0100; 
	if(x==?20'b??1??1?01?0???0?11??) z |= 4'b1000; 
	if(x==?20'b1???????11???0?0?111) z |= 4'b1000; 
	if(x==?20'b????111??1???000???1) z |= 4'b1000; 
	if(x==?20'b????11??110???0??11?) z |= 4'b1000; 
	if(x==?20'b????0?11??11?0??1??1) z |= 4'b0100; 
	if(x==?20'b?1??01?1??11??0??11?) z |= 4'b1100; 
	if(x==?20'b????0?11??11??0?1??1) z |= 4'b0100; 
	if(x==?20'b11???1?011??????1??1) z |= 4'b1000; 
	if(x==?20'b?11??01????10???11??) z |= 4'b0100; 
	if(x==?20'b??11011?????0????11?) z |= 4'b0100; 
	if(x==?20'b??11??1?0?11????1??1) z |= 4'b0100; 
	if(x==?20'b11???110???????0?11?) z |= 4'b1000; 
	if(x==?20'b?1?1??11???10????11?) z |= 4'b0100; 
	if(x==?20'b1?1?11??1??????011??) z |= 4'b1000; 
	if(x==?20'b1????11011???????11?) z |= 4'b1000; 
	if(x==?20'b1???1110?1??????11??) z |= 4'b1000; 
	if(x==?20'b????11??11????001??1) z |= 4'b1000; 
	if(x==?20'b?1???1?01????10?11??) z |= 4'b1000; 
	if(x==?20'b?1?????011?0????1?11) z |= 4'b1000; 
	if(x==?20'b111????011???????1?1) z |= 4'b1000; 
	if(x==?20'b?????111??1?000????1) z |= 4'b0100; 
	if(x==?20'b1???11??1??1?0??1??1) z |= 4'b1000; 
	if(x==?20'b1???11??1??1??0?1??1) z |= 4'b1000; 
	if(x==?20'b11??11??1??????01?1?) z |= 4'b1000; 
	if(x==?20'b1?1??11??11???1??1??) z |= 4'b1000; 
	if(x==?20'b??110?1???11????1??1) z |= 4'b0100; 
	if(x==?20'b???1??????110?0??111) z |= 4'b0100; 
	if(x==?20'b???10111??1?????11??) z |= 4'b0100; 
	if(x==?20'b?1?1??11?0???0??1??1) z |= 4'b0100; 
	if(x==?20'b??1?0???0?11????1?11) z |= 4'b0100; 
	if(x==?20'b?1?1??11?0????0?1??1) z |= 4'b0100; 
	if(x==?20'b??????11?011?0???11?) z |= 4'b0100; 
	if(x==?20'b11??1?10?1???????11?) z |= 4'b1000; 
	if(x==?20'b???1011???11?????11?) z |= 4'b0100; 
	if(x==?20'b11??1??01???????1?11) z |= 4'b1000; 
	if(x==?20'b????11??11???01??11?) z |= 4'b1000; 
	if(x==?20'b??????11??1100??1??1) z |= 4'b0100; 
	if(x==?20'b??11???1?0?1????1?11) z |= 4'b0100; 
	if(x==?20'b?1110?????11?????1?1) z |= 4'b0100; 
	if(x==?20'b??11??11???10???1?1?) z |= 4'b0100; 
	if(x==?20'b?1?1??1101??????11??) z |= 4'b0100; 
	if(x==?20'b11???1??11?????01??1) z |= 4'b1000; 
	if(x==?20'b??11?1?101??????11??) z |= 4'b0100; 
	if(x==?20'b??????11??11?10??11?) z |= 4'b0100; 
	if(x==?20'b1?1?11?0?????0??1??1) z |= 4'b1000; 
	if(x==?20'b?1??1???1?????10111?) z |= 4'b1000; 
	if(x==?20'b1?1?11?0??????0?1??1) z |= 4'b1000; 
	if(x==?20'b1?1?1?1??????0?0?1?1) z |= 4'b1000; 
	if(x==?20'b??1?0?1????1?01?11??) z |= 4'b0100; 
	if(x==?20'b?1?10?11?????0??1??1) z |= 4'b0100; 
	if(x==?20'b?1??0?1????1?01?11??) z |= 4'b0100; 
	if(x==?20'b?1??011??0?1????1??1) z |= 4'b0100; 
	if(x==?20'b11??1?1???10????11??) z |= 4'b1000; 
	if(x==?20'b?1?10?11??????0?1??1) z |= 4'b0100; 
	if(x==?20'b?????11??11??11?1???) z |= 4'b0011; 
	if(x==?20'b11??11??1?1??0???1??) z |= 4'b1000; 
	if(x==?20'b?11?11??110??????1??) z |= 4'b1000; 
	if(x==?20'b11??1??0???1????1?11) z |= 4'b1000; 
	if(x==?20'b??1101?1??1??????11?) z |= 4'b0100; 
	if(x==?20'b11??11??1?1???0??1??) z |= 4'b1000; 
	if(x==?20'b11??11???1?0????1?1?) z |= 4'b1000; 
	if(x==?20'b??110??1???1????1?11) z |= 4'b0100; 
	if(x==?20'b?1??111?1?????00???1) z |= 4'b1000; 
	if(x==?20'b?1?1?1?1????0?0??1?1) z |= 4'b0100; 
	if(x==?20'b??1?111??????1?01??1) z |= 4'b1000; 
	if(x==?20'b?111????00??????1?11) z |= 4'b0100; 
	if(x==?20'b111???????00????1?11) z |= 4'b1000; 
	if(x==?20'b??11??110?1?????1?1?) z |= 4'b0100; 
	if(x==?20'b??11??1???110???1??1) z |= 4'b0100; 
	if(x==?20'b??1??1?0?10???0??11?) z |= 4'b1000; 
	if(x==?20'b??11??11?1?1??0??1??) z |= 4'b0100; 
	if(x==?20'b?11??11?01???1???1??) z |= 4'b0100; 
	if(x==?20'b????11?0??????001?11) z |= 4'b1000; 
	if(x==?20'b111??10?1???????11??) z |= 4'b1000; 
	if(x==?20'b1?1??1??11????1??11?) z |= 4'b1000; 
	if(x==?20'b??1????1???10?1?111?) z |= 4'b0100; 
	if(x==?20'b?1?1??1???11?1???11?) z |= 4'b0100; 
	if(x==?20'b11??1????????0?1111?) z |= 4'b1000; 
	if(x==?20'b11??11?0?1??????1?1?) z |= 4'b1000; 
	if(x==?20'b?1?1??1?01?1????11??) z |= 4'b0100; 
	if(x==?20'b????11??1?1??0?0?11?) z |= 4'b1000; 
	if(x==?20'b??11??11??11?0???1??) z |= 4'b0100; 
	if(x==?20'b????11??1????0001??1) z |= 4'b1000; 
	if(x==?20'b11??1?1??1?????0?11?) z |= 4'b1000; 
	if(x==?20'b1???111??1???00????1) z |= 4'b1000; 
	if(x==?20'b?1??0?1??01??0???11?) z |= 4'b0100; 
	if(x==?20'b??1??111???100?????1) z |= 4'b0100; 
	if(x==?20'b?1???11?1????1?01??1) z |= 4'b1000; 
	if(x==?20'b?111?01????1????11??) z |= 4'b0100; 
	if(x==?20'b??110?11??1?????1?1?) z |= 4'b0100; 
	if(x==?20'b11??1?1????0??0??11?) z |= 4'b1000; 
	if(x==?20'b111??1???10??0???1??) z |= 4'b1000; 
	if(x==?20'b1?1?11?????0?0???11?) z |= 4'b1000; 
	if(x==?20'b?1?1??110?????0??11?) z |= 4'b0100; 
	if(x==?20'b??11?1?10????0???11?) z |= 4'b0100; 
	if(x==?20'b??????11?1?10?0??11?) z |= 4'b0100; 
	if(x==?20'b1?1?11????????001??1) z |= 4'b1000; 
	if(x==?20'b??1?11??1??1???01??1) z |= 4'b1000; 
	if(x==?20'b?1?1??11????00??1??1) z |= 4'b0100; 
	if(x==?20'b?11???11?011?????1??) z |= 4'b0100; 
	if(x==?20'b????11??1????0?11?11) z |= 4'b1000; 
	if(x==?20'b?1???1101??0?????11?) z |= 4'b1000; 
	if(x==?20'b???1?111??1??00????1) z |= 4'b0100; 
	if(x==?20'b??11?1?1??1?0????11?) z |= 4'b0100; 
	if(x==?20'b??????11???1000?1??1) z |= 4'b0100; 
	if(x==?20'b?1???111????0?1?1??1) z |= 4'b0100; 
	if(x==?20'b?1?????01????0?0?111) z |= 4'b1000; 
	if(x==?20'b?111??1??01??0???1??) z |= 4'b0100; 
	if(x==?20'b1?1?1???11???0???1?1) z |= 4'b1000; 
	if(x==?20'b111??1???1?0??0??1??) z |= 4'b1000; 
	if(x==?20'b?111??1??01???0??1??) z |= 4'b0100; 
	if(x==?20'b1????1?011??????1?11) z |= 4'b1000; 
	if(x==?20'b??1?011?0??1?????11?) z |= 4'b0100; 
	if(x==?20'b1?1??1??1??0?0???11?) z |= 4'b1000; 
	if(x==?20'b????111?1??0??0???11) z |= 4'b1000; 
	if(x==?20'b1?1??1??1??0??0??11?) z |= 4'b1000; 
	if(x==?20'b????11?????1?0?11?11) z |= 4'b1000; 
	if(x==?20'b?11??11???10??1??1??) z |= 4'b1000; 
	if(x==?20'b??11??1?????0?1?1?11) z |= 4'b0100; 
	if(x==?20'b?1?1??1?0??1?0???11?) z |= 4'b0100; 
	if(x==?20'b??1??101?1????0??11?) z |= 4'b1000; 
	if(x==?20'b??1?0??????10?0??111) z |= 4'b0100; 
	if(x==?20'b?1?1??1?0??1??0??11?) z |= 4'b0100; 
	if(x==?20'b1?1?111????0??????11) z |= 4'b1000; 
	if(x==?20'b?1?1?1110?????????11) z |= 4'b0100; 
	if(x==?20'b?????1110??1?0????11) z |= 4'b0100; 
	if(x==?20'b??1?11?011??????1??1) z |= 4'b1000; 
	if(x==?20'b??1??11????10?1?1??1) z |= 4'b0100; 
	if(x==?20'b???10?1???11????1?11) z |= 4'b0100; 
	if(x==?20'b????11?0?1???00?1??1) z |= 4'b1000; 
	if(x==?20'b???1011?????0???111?) z |= 4'b0100; 
	if(x==?20'b1????110???????0111?) z |= 4'b1000; 
	if(x==?20'b?11?11??1?1????0?1??) z |= 4'b1000; 
	if(x==?20'b?1?1???1??11??0??1?1) z |= 4'b0100; 
	if(x==?20'b?1???11?1110?????1??) z |= 4'b1000; 
	if(x==?20'b????0?11??1??00?1??1) z |= 4'b0100; 
	if(x==?20'b11??111?1?????0????1) z |= 4'b1000; 
	if(x==?20'b?11???11?1?10????1??) z |= 4'b0100; 
	if(x==?20'b1???1?1?11????0??11?) z |= 4'b1000; 
	if(x==?20'b?1???1101??????0?11?) z |= 4'b1000; 
	if(x==?20'b??1??11?0111?????1??) z |= 4'b0100; 
	if(x==?20'b?1??111??1???0?0???1) z |= 4'b1000; 
	if(x==?20'b1?1?111?11???????1??) z |= 4'b1000; 
	if(x==?20'b??1?111??1????00???1) z |= 4'b1000; 
	if(x==?20'b1???11??1????00?1??1) z |= 4'b1000; 
	if(x==?20'b?1??0?11??11????1??1) z |= 4'b0100; 
	if(x==?20'b????0?1?1???00??111?) z |= 4'b0100; 
	if(x==?20'b1?1???1??1???0?0?1?1) z |= 4'b1000; 
	if(x==?20'b?1??111????0?00????1) z |= 4'b1000; 
	if(x==?20'b??1??1110????00????1) z |= 4'b0100; 
	if(x==?20'b??11?111???1?0?????1) z |= 4'b0100; 
	if(x==?20'b1????110?1???0???11?) z |= 4'b1000; 
	if(x==?20'b?111??110?????????11) z |= 4'b0100; 
	if(x==?20'b??1?011????10????11?) z |= 4'b0100; 
	if(x==?20'b?11???11011??????1??) z |= 4'b0100; 
	if(x==?20'b111?11?????0??????11) z |= 4'b1000; 
	if(x==?20'b????11???1???0001??1) z |= 4'b1000; 
	if(x==?20'b?11?11???110?????1??) z |= 4'b1000; 
	if(x==?20'b?1???111??1?00?????1) z |= 4'b0100; 
	if(x==?20'b?1???1101??????011??) z |= 4'b1000; 
	if(x==?20'b??1??111??1?0?0????1) z |= 4'b0100; 
	if(x==?20'b1?1?11??1??1????1??1) z |= 4'b1000; 
	if(x==?20'b??1?1?1?110?????11??) z |= 4'b1000; 
	if(x==?20'b1?1??1101???????1??1) z |= 4'b1000; 
	if(x==?20'b?1?1011?1???????1??1) z |= 4'b0100; 
	if(x==?20'b?1??1??????0?0?0111?) z |= 4'b1000; 
	if(x==?20'b?1???11??1???1?01??1) z |= 4'b1000; 
	if(x==?20'b??1????10???0?0?111?) z |= 4'b0100; 
	if(x==?20'b???1011???1???0??11?) z |= 4'b0100; 
	if(x==?20'b?1??1?1011???????11?) z |= 4'b1000; 
	if(x==?20'b???1??11???1?00?1??1) z |= 4'b0100; 
	if(x==?20'b?1?1?1????1?0?0??1?1) z |= 4'b0100; 
	if(x==?20'b???1?1?1??11?0???11?) z |= 4'b0100; 
	if(x==?20'b??????11??1?000?1??1) z |= 4'b0100; 
	if(x==?20'b111?11?0??????????11) z |= 4'b1000; 
	if(x==?20'b????111?1?????001??1) z |= 4'b1000; 
	if(x==?20'b?1??11?1??10????11??) z |= 4'b1000; 
	if(x==?20'b?1110?11??????????11) z |= 4'b0100; 
	if(x==?20'b111??1??1??0??????11) z |= 4'b1000; 
	if(x==?20'b11??111?11??????1???) z |= 4'b1000; 
	if(x==?20'b?1?1?111??11?????1??) z |= 4'b0100; 
	if(x==?20'b??1?011????10???11??) z |= 4'b0100; 
	if(x==?20'b?11?1?????00????1?11) z |= 4'b1000; 
	if(x==?20'b??1?11?01????0??1??1) z |= 4'b1000; 
	if(x==?20'b??1????0?1???0?0?111) z |= 4'b1000; 
	if(x==?20'b1???11????????001?11) z |= 4'b1000; 
	if(x==?20'b?1????11?0?1?0??1??1) z |= 4'b0100; 
	if(x==?20'b??1?11?01?????0?1??1) z |= 4'b1000; 
	if(x==?20'b1?1??110???1????1??1) z |= 4'b1000; 
	if(x==?20'b??1?1?1?1????0?0?1?1) z |= 4'b1000; 
	if(x==?20'b?1?1011????1????1??1) z |= 4'b0100; 
	if(x==?20'b?1????11?0?1??0?1??1) z |= 4'b0100; 
	if(x==?20'b?11????100??????1?11) z |= 4'b0100; 
	if(x==?20'b?111??1?0??1??????11) z |= 4'b0100; 
	if(x==?20'b1?1?111????0?????11?) z |= 4'b1000; 
	if(x==?20'b?1?1?1110????????11?) z |= 4'b0100; 
	if(x==?20'b1?1?1????????0?0?111) z |= 4'b1000; 
	if(x==?20'b?1??11??11?0????1?1?) z |= 4'b1000; 
	if(x==?20'b?1??0?????1?0?0??111) z |= 4'b0100; 
	if(x==?20'b?11?0110?????0???11?) z |= 4'b1100; 
	if(x==?20'b?1?1???1????0?0??111) z |= 4'b0100; 
	if(x==?20'b?11?0110??????0??11?) z |= 4'b1100; 
	if(x==?20'b?11?1?1??10???0??1??) z |= 4'b1000; 
	if(x==?20'b?1??0?11???1?0??1??1) z |= 4'b0100; 
	if(x==?20'b111?11??1?1??????1??) z |= 4'b1000; 
	if(x==?20'b??1??11???1?0?1?1??1) z |= 4'b0100; 
	if(x==?20'b?1??011?0?1?????11??) z |= 4'b0100; 
	if(x==?20'b?1?1??1???1??10??11?) z |= 4'b0100; 
	if(x==?20'b?1??0?11???1??0?1??1) z |= 4'b0100; 
	if(x==?20'b??1?01?1??11?????11?) z |= 4'b0100; 
	if(x==?20'b?1??1???1????0?1111?) z |= 4'b1000; 
	if(x==?20'b?1??11?011??????1?1?) z |= 4'b1000; 
	if(x==?20'b?1???1?1?011????11??) z |= 4'b0100; 
	if(x==?20'b11??????1????0?0?111) z |= 4'b1000; 
	if(x==?20'b?1??111??????000???1) z |= 4'b1000; 
	if(x==?20'b?1??1?1?11?????0?11?) z |= 4'b1000; 
	if(x==?20'b????111?11???00????1) z |= 4'b1000; 
	if(x==?20'b111??110?1???????1??) z |= 4'b1000; 
	if(x==?20'b??11?111??11????1???) z |= 4'b0100; 
	if(x==?20'b?1???1?1???10?0??1?1) z |= 4'b0100; 
	if(x==?20'b1???1?10??????0?111?) z |= 4'b1000; 
	if(x==?20'b?111??11?1?1?????1??) z |= 4'b0100; 
	if(x==?20'b?1??1????10??00?11??) z |= 4'b1000; 
	if(x==?20'b?11?????00?1????1?11) z |= 4'b0100; 
	if(x==?20'b??1??111????000????1) z |= 4'b0100; 
	if(x==?20'b??1???110?11????1?1?) z |= 4'b0100; 
	if(x==?20'b1?1??1???1???01??11?) z |= 4'b1000; 
	if(x==?20'b?1??1?1?1??0??0??11?) z |= 4'b1000; 
	if(x==?20'b11???1101????????11?) z |= 4'b1000; 
	if(x==?20'b?11??1??110??0???1??) z |= 4'b1000; 
	if(x==?20'b111?1??????????1111?) z |= 4'b1000; 
	if(x==?20'b???101?1?????0??111?) z |= 4'b0100; 
	if(x==?20'b?111011???1??????1??) z |= 4'b0100; 
	if(x==?20'b??1?11??1?????001??1) z |= 4'b1000; 
	if(x==?20'b?11??1?1?01??0???1??) z |= 4'b0100; 
	if(x==?20'b1?1?111??1????0????1) z |= 4'b1000; 
	if(x==?20'b??11???????10?0??111) z |= 4'b0100; 
	if(x==?20'b??1?11??1?0??0??11??) z |= 4'b1000; 
	if(x==?20'b1?1?????1????0?011?1) z |= 4'b1000; 
	if(x==?20'b?11??1??001?????11??) z |= 4'b0100; 
	if(x==?20'b??1??110?1?????0?11?) z |= 4'b1000; 
	if(x==?20'b?1????11????0?1?1?11) z |= 4'b0100; 
	if(x==?20'b?1??1?101?????0??11?) z |= 4'b1000; 
	if(x==?20'b?11??1??11?0??0??1??) z |= 4'b1000; 
	if(x==?20'b?1???01?????0?0?111?) z |= 4'b0100; 
	if(x==?20'b??1?011?0?????0??11?) z |= 4'b0100; 
	if(x==?20'b??1?0?11??11????1?1?) z |= 4'b0100; 
	if(x==?20'b??1??10??????0?0111?) z |= 4'b1000; 
	if(x==?20'b??11011????1?????11?) z |= 4'b0100; 
	if(x==?20'b??1????1?01??00?11??) z |= 4'b0100; 
	if(x==?20'b??1??1?10??1?0???11?) z |= 4'b0100; 
	if(x==?20'b1???11???1???00?1??1) z |= 4'b1000; 
	if(x==?20'b?1?1?111??1??0?????1) z |= 4'b0100; 
	if(x==?20'b?1???110???0?0???11?) z |= 4'b1000; 
	if(x==?20'b?1??011???1?0????11?) z |= 4'b0100; 
	if(x==?20'b?1????11???100??1??1) z |= 4'b0100; 
	if(x==?20'b?????111??11?00????1) z |= 4'b0100; 
	if(x==?20'b??1??1?1??110????11?) z |= 4'b0100; 
	if(x==?20'b?1?1???10????0??111?) z |= 4'b0100; 
	if(x==?20'b??1?111??????0?11??1) z |= 4'b1000; 
	if(x==?20'b??1?1???11?0????1?11) z |= 4'b1000; 
	if(x==?20'b1?1?1??????0??0?111?) z |= 4'b1000; 
	if(x==?20'b?1??1???11?0????1?11) z |= 4'b1000; 
	if(x==?20'b?11???1??011?0???1??) z |= 4'b0100; 
	if(x==?20'b?1?1???????10?0?11?1) z |= 4'b0100; 
	if(x==?20'b??1?111?1??0??????11) z |= 4'b1000; 
	if(x==?20'b???1??11??1??00?1??1) z |= 4'b0100; 
	if(x==?20'b?11???1??011??0??1??) z |= 4'b0100; 
	if(x==?20'b????111????0?00???11) z |= 4'b1000; 
	if(x==?20'b?????1110????00???11) z |= 4'b0100; 
	if(x==?20'b??1?01?1???1?0???11?) z |= 4'b0100; 
	if(x==?20'b??11???1?????10?111?) z |= 4'b0100; 
	if(x==?20'b?????1101??????0111?) z |= 4'b1000; 
	if(x==?20'b?1??1??011??????1?11) z |= 4'b1000; 
	if(x==?20'b1???111?11??????11??) z |= 4'b1000; 
	if(x==?20'b????111??1????001??1) z |= 4'b1000; 
	if(x==?20'b?1???1110??1??????11) z |= 4'b0100; 
	if(x==?20'b??1?11?0?1???0??1??1) z |= 4'b1000; 
	if(x==?20'b11???1???????0?11?11) z |= 4'b1000; 
	if(x==?20'b??1?11?0?1????0?1??1) z |= 4'b1000; 
	if(x==?20'b??1????10?11????1?11) z |= 4'b0100; 
	if(x==?20'b?1?????10?11????1?11) z |= 4'b0100; 
	if(x==?20'b????011????10???111?) z |= 4'b0100; 
	if(x==?20'b?1??0?11??1??0??1??1) z |= 4'b0100; 
	if(x==?20'b111?111?1??????????1) z |= 4'b1000; 
	if(x==?20'b?1??1?10???????0111?) z |= 4'b1000; 
	if(x==?20'b11??111??????00????1) z |= 4'b1000; 
	if(x==?20'b11??1?1?11???????11?) z |= 4'b1000; 
	if(x==?20'b?1??0?11??1???0?1??1) z |= 4'b0100; 
	if(x==?20'b111??1?01???????11??) z |= 4'b1000; 
	if(x==?20'b??1???11011?????1?1?) z |= 4'b0100; 
	if(x==?20'b?1??11???110????1?1?) z |= 4'b1000; 
	if(x==?20'b??11?111?????00????1) z |= 4'b0100; 
	if(x==?20'b??1?0??1??11????1?11) z |= 4'b0100; 
	if(x==?20'b??1?01?1????0???111?) z |= 4'b0100; 
	if(x==?20'b?????11011???0???11?) z |= 4'b1000; 
	if(x==?20'b?????11011????0??11?) z |= 4'b1000; 
	if(x==?20'b???1?111??11????11??) z |= 4'b0100; 
	if(x==?20'b1?1?11??1????0??1??1) z |= 4'b1000; 
	if(x==?20'b?11????011???0???1?1) z |= 4'b1000; 
	if(x==?20'b1?1?11??1?????0?1??1) z |= 4'b1000; 
	if(x==?20'b?1110?1????1????11??) z |= 4'b0100; 
	if(x==?20'b?11????011????0??1?1) z |= 4'b1000; 
	if(x==?20'b??11??1?????000??11?) z |= 4'b0100; 
	if(x==?20'b11??1???1??1????1?11) z |= 4'b1000; 
	if(x==?20'b11???1???????000?11?) z |= 4'b1000; 
	if(x==?20'b?111?111???1???????1) z |= 4'b0100; 
	if(x==?20'b1?1??110?1???????11?) z |= 4'b1000; 
	if(x==?20'b??1?11???1????001??1) z |= 4'b1000; 
	if(x==?20'b1?1?11?????1?0??1??1) z |= 4'b1000; 
	if(x==?20'b?11?1111?11??????1??) z |= 4'b1100; 
	if(x==?20'b1?1?11?????1??0?1??1) z |= 4'b1000; 
	if(x==?20'b?1?1011???1??????11?) z |= 4'b0100; 
	if(x==?20'b?1?1??11???1?0??1??1) z |= 4'b0100; 
	if(x==?20'b????11??1?????001?11) z |= 4'b1000; 
	if(x==?20'b?1??1?10?1???0???11?) z |= 4'b1000; 
	if(x==?20'b????011???11?0???11?) z |= 4'b0100; 
	if(x==?20'b?1?1??11???1??0?1??1) z |= 4'b0100; 
	if(x==?20'b?11???1?011??0???1??) z |= 4'b0100; 
	if(x==?20'b??1?1?10?1????0??11?) z |= 4'b1000; 
	if(x==?20'b??11?1?1??11?????11?) z |= 4'b0100; 
	if(x==?20'b11??11??11??????1?1?) z |= 4'b1000; 
	if(x==?20'b?1????11??1?00??1??1) z |= 4'b0100; 
	if(x==?20'b?111???1?0??????1?11) z |= 4'b0100; 
	if(x==?20'b????011???11??0??11?) z |= 4'b0100; 
	if(x==?20'b?11?0?????11?0???1?1) z |= 4'b0100; 
	if(x==?20'b????111??????0001??1) z |= 4'b1000; 
	if(x==?20'b111??1??1??????011??) z |= 4'b1000; 
	if(x==?20'b?11?0?????11??0??1?1) z |= 4'b0100; 
	if(x==?20'b?1????11??1??10??11?) z |= 4'b0100; 
	if(x==?20'b??11011??1??????11??) z |= 4'b0100; 
	if(x==?20'b?11??1???110??0??1??) z |= 4'b1000; 
	if(x==?20'b?????111????000?1??1) z |= 4'b0100; 
	if(x==?20'b111?1??0????????1?11) z |= 4'b1000; 
	if(x==?20'b????11?????1??001?11) z |= 4'b1000; 
	if(x==?20'b??1?11???1???01??11?) z |= 4'b1000; 
	if(x==?20'b1????1101???????111?) z |= 4'b1000; 
	if(x==?20'b?1??01?1??1??0???11?) z |= 4'b0100; 
	if(x==?20'b11???110??1?????11??) z |= 4'b1000; 
	if(x==?20'b?111??1????10???11??) z |= 4'b0100; 
	if(x==?20'b??1?01?1??1???0??11?) z |= 4'b0100; 
	if(x==?20'b?1110??1????????1?11) z |= 4'b0100; 
	if(x==?20'b111?11???1???0???1??) z |= 4'b1000; 
	if(x==?20'b??1?111?1??0????11??) z |= 4'b1000; 
	if(x==?20'b111?11???1????0??1??) z |= 4'b1000; 
	if(x==?20'b?11?1?????????10111?) z |= 4'b1000; 
	if(x==?20'b?11??11011???????1??) z |= 4'b1000; 
	if(x==?20'b11??1?1?1?????0??11?) z |= 4'b1000; 
	if(x==?20'b1?1?11??1????0???11?) z |= 4'b1000; 
	if(x==?20'b????1?101?????0?111?) z |= 4'b1000; 
	if(x==?20'b?11????1????0?1?111?) z |= 4'b0100; 
	if(x==?20'b??11??11??11????1?1?) z |= 4'b0100; 
	if(x==?20'b???1011????1????111?) z |= 4'b0100; 
	if(x==?20'b??1??1??11???01??11?) z |= 4'b1000; 
	if(x==?20'b?111??11??1??0???1??) z |= 4'b0100; 
	if(x==?20'b?1????1???11?10??11?) z |= 4'b0100; 
	if(x==?20'b?11??1101?1??????1??) z |= 4'b1000; 
	if(x==?20'b?111??11??1???0??1??) z |= 4'b0100; 
	if(x==?20'b?1??1?1??1???0?0?11?) z |= 4'b1000; 
	if(x==?20'b?11?111???????00???1) z |= 4'b1000; 
	if(x==?20'b??1?111?11????0????1) z |= 4'b1000; 
	if(x==?20'b??1?11???1???0?0?11?) z |= 4'b1000; 
	if(x==?20'b11??1?10????????111?) z |= 4'b1000; 
	if(x==?20'b111??1??11????0??1??) z |= 4'b1000; 
	if(x==?20'b?1???111?0?1????11??) z |= 4'b0100; 
	if(x==?20'b?11??111????00?????1) z |= 4'b0100; 
	if(x==?20'b?11?011??1?1?????1??) z |= 4'b0100; 
	if(x==?20'b11???110?????0???11?) z |= 4'b1000; 
	if(x==?20'b??11011??????0???11?) z |= 4'b0100; 
	if(x==?20'b??1?1???1?0???0?111?) z |= 4'b1000; 
	if(x==?20'b??1101?1????????111?) z |= 4'b0100; 
	if(x==?20'b11???110??????0??11?) z |= 4'b1000; 
	if(x==?20'b??11011???????0??11?) z |= 4'b0100; 
	if(x==?20'b??1?11???????0001??1) z |= 4'b1000; 
	if(x==?20'b?1?1??11???1??0??11?) z |= 4'b0100; 
	if(x==?20'b??11?1?1???1?0???11?) z |= 4'b0100; 
	if(x==?20'b?11?1??11??1????1?11) z |= 4'b1100; 
	if(x==?20'b????01?1???1?0??111?) z |= 4'b0100; 
	if(x==?20'b????11??11???00?1??1) z |= 4'b1000; 
	if(x==?20'b?11?011???11?????1??) z |= 4'b0100; 
	if(x==?20'b?1????11????000?1??1) z |= 4'b0100; 
	if(x==?20'b?111????111???????11) z |= 4'b0100; 
	if(x==?20'b?1????11??1?0?0??11?) z |= 4'b0100; 
	if(x==?20'b??1??1?1??1?0?0??11?) z |= 4'b0100; 
	if(x==?20'b11??111?1?????????11) z |= 4'b1000; 
	if(x==?20'b11??11??1????0??1?1?) z |= 4'b1000; 
	if(x==?20'b?111??1???11?0???1??) z |= 4'b0100; 
	if(x==?20'b11??11??1?????0?1?1?) z |= 4'b1000; 
	if(x==?20'b111??????111??????11) z |= 4'b1000; 
	if(x==?20'b?1???111??11?0?????1) z |= 4'b0100; 
	if(x==?20'b?11????0?????0?0?111) z |= 4'b1000; 
	if(x==?20'b?1?1??11???1??0?11??) z |= 4'b0100; 
	if(x==?20'b?11?0???????0?0??111) z |= 4'b0100; 
	if(x==?20'b??1?111??0???0????11) z |= 4'b0100; 
	if(x==?20'b?1???111??0???0???11) z |= 4'b1000; 
	if(x==?20'b?1?????1?0?1?0??111?) z |= 4'b0100; 
	if(x==?20'b?1???1110????0????11) z |= 4'b0100; 
	if(x==?20'b??1?111????0??0???11) z |= 4'b1000; 
	if(x==?20'b??11??11???1?0??1?1?) z |= 4'b0100; 
	if(x==?20'b??11?111???1??????11) z |= 4'b0100; 
	if(x==?20'b11???1??11???0??1??1) z |= 4'b1000; 
	if(x==?20'b?11??11?????0?1?1??1) z |= 4'b0100; 
	if(x==?20'b??????11??11?00?1??1) z |= 4'b0100; 
	if(x==?20'b??11??11???1??0?1?1?) z |= 4'b0100; 
	if(x==?20'b11???1??11????0?1??1) z |= 4'b1000; 
	if(x==?20'b?????111111???????11) z |= 4'b1000; 
	if(x==?20'b?11??11?11?0????1?1?) z |= 4'b1100; 
	if(x==?20'b??1????1???1?10?111?) z |= 4'b0100; 
	if(x==?20'b????111??111??????11) z |= 4'b0100; 
	if(x==?20'b?1??111?1????00????1) z |= 4'b1000; 
	if(x==?20'b?11??11011??????1?1?) z |= 4'b1100; 
	if(x==?20'b?1??11???????000?11?) z |= 4'b1000; 
	if(x==?20'b?11??1??11?0????1??1) z |= 4'b1000; 
	if(x==?20'b111?11??1?????????11) z |= 4'b1000; 
	if(x==?20'b??1???11????000??11?) z |= 4'b0100; 
	if(x==?20'b??11??1???11?0??1??1) z |= 4'b0100; 
	if(x==?20'b?11??11?0?11????1?1?) z |= 4'b1100; 
	if(x==?20'b?111???1??????1?111?) z |= 4'b0100; 
	if(x==?20'b??11??1???11??0?1??1) z |= 4'b0100; 
	if(x==?20'b????0?11?????00?1?11) z |= 4'b0100; 
	if(x==?20'b??1?????11???0?0?111) z |= 4'b1000; 
	if(x==?20'b11??1?1??1???0???11?) z |= 4'b1000; 
	if(x==?20'b1?1??11?1??1????1??1) z |= 4'b1000; 
	if(x==?20'b111?111???????0????1) z |= 4'b1000; 
	if(x==?20'b?1?1?11?1??1????1??1) z |= 4'b0100; 
	if(x==?20'b1?1?1?1??1????0??11?) z |= 4'b1000; 
	if(x==?20'b?11??1?011??????1??1) z |= 4'b1000; 
	if(x==?20'b?111?111?????0?????1) z |= 4'b0100; 
	if(x==?20'b?11?011?????0????11?) z |= 4'b0100; 
	if(x==?20'b?11??110???????0?11?) z |= 4'b1000; 
	if(x==?20'b?11???1?0?11????1??1) z |= 4'b0100; 
	if(x==?20'b?1???1??1????000?11?) z |= 4'b1000; 
	if(x==?20'b??1??11011???????11?) z |= 4'b1000; 
	if(x==?20'b??1??111???1?00????1) z |= 4'b0100; 
	if(x==?20'b1?1??1?1?1????0??11?) z |= 4'b1000; 
	if(x==?20'b?111??11???1??????11) z |= 4'b0100; 
	if(x==?20'b?11?011???11????1?1?) z |= 4'b1100; 
	if(x==?20'b1?1?11???????00?1??1) z |= 4'b1000; 
	if(x==?20'b??1?11??1??1?0??1??1) z |= 4'b1000; 
	if(x==?20'b?1??11??111???????11) z |= 4'b1000; 
	if(x==?20'b??????1?001?1???11??) z |= 4'b0100; 
	if(x==?20'b??1?11??1??1??0?1??1) z |= 4'b1000; 
	if(x==?20'b1?1?111?1????????11?) z |= 4'b1000; 
	if(x==?20'b?1?1??11?????00?1??1) z |= 4'b0100; 
	if(x==?20'b?1?1?1?1??1??0???11?) z |= 4'b0100; 
	if(x==?20'b??1?01??????00??111?) z |= 4'b0100; 
	if(x==?20'b?1??111???????00??11) z |= 4'b1000; 
	if(x==?20'b?1????10??????00111?) z |= 4'b1000; 
	if(x==?20'b?11?11??1??????01?1?) z |= 4'b1000; 
	if(x==?20'b??1???1????1000??11?) z |= 4'b0100; 
	if(x==?20'b??11?1?1??1???0??11?) z |= 4'b0100; 
	if(x==?20'b111?111??1????????1?) z |= 4'b1000; 
	if(x==?20'b??1??111????00????11) z |= 4'b0100; 
	if(x==?20'b?11?0?1???11????1??1) z |= 4'b0100; 
	if(x==?20'b?1????????110?0??111) z |= 4'b0100; 
	if(x==?20'b?????1???100???111??) z |= 4'b1000; 
	if(x==?20'b????11???????0001?11) z |= 4'b1000; 
	if(x==?20'b?11?1?10?1???????11?) z |= 4'b1000; 
	if(x==?20'b??1???11?111??????11) z |= 4'b0100; 
	if(x==?20'b?1??011???11?????11?) z |= 4'b0100; 
	if(x==?20'b?11?1??01???????1?11) z |= 4'b1000; 
	if(x==?20'b??????11????000?1?11) z |= 4'b0100; 
	if(x==?20'b111??11?1?1??????1??) z |= 4'b1000; 
	if(x==?20'b?111?111??1???????1?) z |= 4'b0100; 
	if(x==?20'b?11???11???10???1?1?) z |= 4'b0100; 
	if(x==?20'b?1?1?111???1?????11?) z |= 4'b0100; 
	if(x==?20'b?11??1??11?????01??1) z |= 4'b1000; 
	if(x==?20'b?11??1?101??????11??) z |= 4'b0100; 
	if(x==?20'b????111?111???????1?) z |= 4'b0010; 
	if(x==?20'b?111?11??1?1?????1??) z |= 4'b0100; 
	if(x==?20'b1????110?????0??111?) z |= 4'b1000; 
	if(x==?20'b11??111?1???????1?1?) z |= 4'b1000; 
	if(x==?20'b?11?1?1???10????11??) z |= 4'b1000; 
	if(x==?20'b?11?11??1?1??0???1??) z |= 4'b1000; 
	if(x==?20'b?11?1??0???1????1?11) z |= 4'b1000; 
	if(x==?20'b???1011???????0?111?) z |= 4'b0100; 
	if(x==?20'b?11?01?1??1??????11?) z |= 4'b0100; 
	if(x==?20'b?11?11??1?1???0??1??) z |= 4'b1000; 
	if(x==?20'b?11?11???1?0????1?1?) z |= 4'b1000; 
	if(x==?20'b?11?0??1???1????1?11) z |= 4'b0100; 
	if(x==?20'b?1??1?101???????111?) z |= 4'b1000; 
	if(x==?20'b?11???110?1?????1?1?) z |= 4'b0100; 
	if(x==?20'b?11???11?1?1?0???1??) z |= 4'b0100; 
	if(x==?20'b11???1????????001?11) z |= 4'b1000; 
	if(x==?20'b?11???1???110???1??1) z |= 4'b0100; 
	if(x==?20'b?11???11?1?1??0??1??) z |= 4'b0100; 
	if(x==?20'b?????111?111??????1?) z |= 4'b0001; 
	if(x==?20'b?1???1101????0???11?) z |= 4'b1000; 
	if(x==?20'b?11?1????????0?1111?) z |= 4'b1000; 
	if(x==?20'b?11?11?0?1??????1?1?) z |= 4'b1000; 
	if(x==?20'b111??????????0?0?111) z |= 4'b1000; 
	if(x==?20'b?11?1?1??1?????0?11?) z |= 4'b1000; 
	if(x==?20'b??11?111???1????1?1?) z |= 4'b0100; 
	if(x==?20'b??1?111??1???00????1) z |= 4'b1000; 
	if(x==?20'b?111????????0?0??111) z |= 4'b0100; 
	if(x==?20'b????11????00???01??1) z |= 4'b1000; 
	if(x==?20'b??????1100??0???1??1) z |= 4'b0100; 
	if(x==?20'b????0?1?1????00?111?) z |= 4'b0100; 
	if(x==?20'b?11?0?11??1?????1?1?) z |= 4'b0100; 
	if(x==?20'b?11?1?1????0??0??11?) z |= 4'b1000; 
	if(x==?20'b111??110?????????11?) z |= 4'b1000; 
	if(x==?20'b?111011??????????11?) z |= 4'b0100; 
	if(x==?20'b?11??1?10????0???11?) z |= 4'b0100; 
	if(x==?20'b?11??1???????1?01?11) z |= 4'b1000; 
	if(x==?20'b??1?01?1???1????111?) z |= 4'b0100; 
	if(x==?20'b??1?011????1??0??11?) z |= 4'b0100; 
	if(x==?20'b?1???1101????0??11??) z |= 4'b1000; 
	if(x==?20'b?1???111??1??00????1) z |= 4'b0100; 
	if(x==?20'b?11??1?1??1?0????11?) z |= 4'b0100; 
	if(x==?20'b11??111???????0???11) z |= 4'b1000; 
	if(x==?20'b111?11??1???????1?1?) z |= 4'b1000; 
	if(x==?20'b??1??1?011??????1?11) z |= 4'b1000; 
	if(x==?20'b??11?111?????0????11) z |= 4'b0100; 
	if(x==?20'b?11???1?????0?1?1?11) z |= 4'b0100; 
	if(x==?20'b??1?011????1??0?11??) z |= 4'b0100; 
	if(x==?20'b???1??11?????00?1?11) z |= 4'b0100; 
	if(x==?20'b?111??11???1????1?1?) z |= 4'b0100; 
	if(x==?20'b111??1??11??????1??1) z |= 4'b1000; 
	if(x==?20'b111??11????????0?11?) z |= 4'b1000; 
	if(x==?20'b?1??0?1???11????1?11) z |= 4'b0100; 
	if(x==?20'b?111?11?????0????11?) z |= 4'b0100; 
	if(x==?20'b?1??011?????0???111?) z |= 4'b0100; 
	if(x==?20'b??1??110???????0111?) z |= 4'b1000; 
	if(x==?20'b1?1?111??1??????11??) z |= 4'b1000; 
	if(x==?20'b1????10??10?????11??) z |= 4'b1000; 
	if(x==?20'b???11??1?1??1???11??) z |= 4'b0100; 
	if(x==?20'b?????1?0???1?00?111?) z |= 4'b1001; 
	if(x==?20'b11????1???????00111?) z |= 4'b1000; 
	if(x==?20'b?1??1?1?11???0???11?) z |= 4'b1000; 
	if(x==?20'b??11?1??????00??111?) z |= 4'b0100; 
	if(x==?20'b?11?111?1?????0????1) z |= 4'b1000; 
	if(x==?20'b??1?1?1?11????0??11?) z |= 4'b1000; 
	if(x==?20'b???11??1??1?1???11??) z |= 4'b0100; 
	if(x==?20'b???1?01??01?????11??) z |= 4'b0100; 
	if(x==?20'b11??111??1??????1?1?) z |= 4'b1000; 
	if(x==?20'b?11?0??1??1?????1?11) z |= 4'b0100; 
	if(x==?20'b?????1?????1?000111?) z |= 4'b1000; 
	if(x==?20'b111?11????????0???11) z |= 4'b1000; 
	if(x==?20'b?111??1???11????1??1) z |= 4'b0100; 
	if(x==?20'b?1?1?111??1?????11??) z |= 4'b0100; 
	if(x==?20'b?111??11?????0????11) z |= 4'b0100; 
	if(x==?20'b??1??1?111????0??11?) z |= 4'b1000; 
	if(x==?20'b??1?11??1????00?1??1) z |= 4'b1000; 
	if(x==?20'b111?1?1??1???????11?) z |= 4'b1000; 
	if(x==?20'b1???1??1?1?????111??) z |= 4'b1000; 
	if(x==?20'b111?1???1???????1?11) z |= 4'b1000; 
	if(x==?20'b1???11????00????1??1) z |= 4'b1000; 
	if(x==?20'b??????1?1???000?111?) z |= 4'b0110; 
	if(x==?20'b??11?111??1?????1?1?) z |= 4'b0100; 
	if(x==?20'b???1??1100??????1??1) z |= 4'b0100; 
	if(x==?20'b?11??111???1?0?????1) z |= 4'b0100; 
	if(x==?20'b??11?11?11??????1?1?) z |= 4'b0100; 
	if(x==?20'b1???1??1??1????111??) z |= 4'b1000; 
	if(x==?20'b111?1??????1????1?11) z |= 4'b1000; 
	if(x==?20'b?1???110?????00?1??1) z |= 4'b1000; 
	if(x==?20'b??1?011??????00?1??1) z |= 4'b0100; 
	if(x==?20'b?111?1?1??1??????11?) z |= 4'b0100; 
	if(x==?20'b?1????11???1?00?1??1) z |= 4'b0100; 
	if(x==?20'b?1???1?1??11?0???11?) z |= 4'b0100; 
	if(x==?20'b??1??1?1??11??0??11?) z |= 4'b0100; 
	if(x==?20'b?111???1???1????1?11) z |= 4'b0100; 
	if(x==?20'b?11?111?11??????1???) z |= 4'b1000; 
	if(x==?20'b??1?11????????001?11) z |= 4'b1000; 
	if(x==?20'b11???11???11????1?1?) z |= 4'b1000; 
	if(x==?20'b?????1101????0??111?) z |= 4'b1000; 
	if(x==?20'b111?11???1??????1?1?) z |= 4'b1000; 
	if(x==?20'b?111??11??1?????1?1?) z |= 4'b0100; 
	if(x==?20'b1?1??110????????111?) z |= 4'b1000; 
	if(x==?20'b?1?1011?????????111?) z |= 4'b0100; 
	if(x==?20'b????011????1??0?111?) z |= 4'b0100; 
	if(x==?20'b?????1???100?1??11??) z |= 4'b1000; 
	if(x==?20'b?1???11??????0001??1) z |= 4'b1000; 
	if(x==?20'b??1??11?????000?1??1) z |= 4'b0100; 
	if(x==?20'b?11?????1????0?0?111) z |= 4'b1000; 
	if(x==?20'b?1??1?10?????0??111?) z |= 4'b1000; 
	if(x==?20'b?11??111??11????1???) z |= 4'b0100; 
	if(x==?20'b??????1?001??1??11??) z |= 4'b0100; 
	if(x==?20'b??1?1?10??????0?111?) z |= 4'b1000; 
	if(x==?20'b1?1??1??11??????1?11) z |= 4'b1000; 
	if(x==?20'b?1??01?1?????0??111?) z |= 4'b0100; 
	if(x==?20'b??1?01?1??????0?111?) z |= 4'b0100; 
	if(x==?20'b????01101??1?????1?1) z |= 4'b1100; 
	if(x==?20'b?11????????10?0??111) z |= 4'b0100; 
	if(x==?20'b?????1???100??1?11??) z |= 4'b1000; 
	if(x==?20'b?1??111?1?????0???11) z |= 4'b1000; 
	if(x==?20'b?1????101?????0?111?) z |= 4'b1000; 
	if(x==?20'b??????1?001???1?11??) z |= 4'b0100; 
	if(x==?20'b??1?11???1???00?1??1) z |= 4'b1000; 
	if(x==?20'b?1?1??1???11????1?11) z |= 4'b0100; 
	if(x==?20'b?111111???????????11) z |= 4'b0100; 
	if(x==?20'b111??1???1????0???11) z |= 4'b1000; 
	if(x==?20'b??1?01?????1?0??111?) z |= 4'b0100; 
	if(x==?20'b111??111??????????11) z |= 4'b1000; 
	if(x==?20'b?1????11??1??00?1??1) z |= 4'b0100; 
	if(x==?20'b111??1??1????0??11??) z |= 4'b1000; 
	if(x==?20'b??1??111???1?0????11) z |= 4'b0100; 
	if(x==?20'b?111??1???1??0????11) z |= 4'b0100; 
	if(x==?20'b111??1??1?????0?11??) z |= 4'b1000; 
	if(x==?20'b1???111?1?0????????1) z |= 4'b1000; 
	if(x==?20'b?11????1?????10?111?) z |= 4'b0100; 
	if(x==?20'b????1?1??1??1?1??1??) z |= 4'b0010; 
	if(x==?20'b??1?111?11??????11??) z |= 4'b1000; 
	if(x==?20'b??????11???1?00?1?11) z |= 4'b0100; 
	if(x==?20'b?111??1????1?0??11??) z |= 4'b0100; 
	if(x==?20'b?111??1????1??0?11??) z |= 4'b0100; 
	if(x==?20'b?1????1?1?????00111?) z |= 4'b1000; 
	if(x==?20'b?1??111?11??????1?1?) z |= 4'b1000; 
	if(x==?20'b?????1?1??1??1?1?1??) z |= 4'b0001; 
	if(x==?20'b?1?1?11???1??0???11?) z |= 4'b0100; 
	if(x==?20'b11???11??????00?1??1) z |= 4'b1000; 
	if(x==?20'b???1?111?0?1???????1) z |= 4'b0100; 
	if(x==?20'b?11?111??????00????1) z |= 4'b1000; 
	if(x==?20'b??11?11??????00?1??1) z |= 4'b0100; 
	if(x==?20'b?11?1?1?11???????11?) z |= 4'b1000; 
	if(x==?20'b??1??1?????100??111?) z |= 4'b0100; 
	if(x==?20'b????11??1?00????1??1) z |= 4'b1000; 
	if(x==?20'b?11??111?????00????1) z |= 4'b0100; 
	if(x==?20'b?????1??1?1?1?1??1??) z |= 4'b0010; 
	if(x==?20'b??????1??1?1?1?1?1??) z |= 4'b0001; 
	if(x==?20'b?1???111??11????11??) z |= 4'b0100; 
	if(x==?20'b?????1??1?1??1?1?11?) z |= 4'b1000; 
	if(x==?20'b?1???10??10???0??1??) z |= 4'b1000; 
	if(x==?20'b??????1?1?1?1?1??11?) z |= 4'b0100; 
	if(x==?20'b?11???1?????000??11?) z |= 4'b0100; 
	if(x==?20'b?????1???1?1?1?1?11?) z |= 4'b1000; 
	if(x==?20'b??????1??1?11?1??11?) z |= 4'b0100; 
	if(x==?20'b?11??1???????000?11?) z |= 4'b1000; 
	if(x==?20'b??1??01??01??0???1??) z |= 4'b0100; 
	if(x==?20'b????011?00??????1??1) z |= 4'b0100; 
	if(x==?20'b??1??111??11????1?1?) z |= 4'b0100; 
	if(x==?20'b?????110??00????1??1) z |= 4'b1000; 
	if(x==?20'b??????1100?1????1??1) z |= 4'b0100; 
	if(x==?20'b111?1????1??????111?) z |= 4'b1000; 
	if(x==?20'b?11?11??11??????1?1?) z |= 4'b1000; 
	if(x==?20'b?11??1?1??11?????11?) z |= 4'b0100; 
	if(x==?20'b1???1??1?1???1??11??) z |= 4'b1000; 
	if(x==?20'b???11??1?1???1??11??) z |= 4'b0100; 
	if(x==?20'b?111???1??1?????111?) z |= 4'b0100; 
	if(x==?20'b?11?011??1??????11??) z |= 4'b0100; 
	if(x==?20'b??1??1101???????111?) z |= 4'b1000; 
	if(x==?20'b1???1??1??1??1??11??) z |= 4'b1000; 
	if(x==?20'b???11??1??1??1??11??) z |= 4'b0100; 
	if(x==?20'b?11??110??1?????11??) z |= 4'b1000; 
	if(x==?20'b???1?1??1??11???11??) z |= 4'b0100; 
	if(x==?20'b1????1?0?10?????11??) z |= 4'b1000; 
	if(x==?20'b11????1?1?????0?111?) z |= 4'b1000; 
	if(x==?20'b??????11??1??00?1?11) z |= 4'b0100; 
	if(x==?20'b?11?1?1?1?????0??11?) z |= 4'b1000; 
	if(x==?20'b111?111?????????1?1?) z |= 4'b1000; 
	if(x==?20'b1???1??1?1????1?11??) z |= 4'b1000; 
	if(x==?20'b?11???11??11????1?1?) z |= 4'b0100; 
	if(x==?20'b???11??1?1????1?11??) z |= 4'b0100; 
	if(x==?20'b?1??011????1????111?) z |= 4'b0100; 
	if(x==?20'b?111?111????????1?1?) z |= 4'b0100; 
	if(x==?20'b?11??11???????001??1) z |= 4'b1000; 
	if(x==?20'b???10?1??01?????11??) z |= 4'b0100; 
	if(x==?20'b1?????1?1??1???111??) z |= 4'b1000; 
	if(x==?20'b1???1??1??1???1?11??) z |= 4'b1000; 
	if(x==?20'b?11?1?10????????111?) z |= 4'b1000; 
	if(x==?20'b???11??1??1???1?11??) z |= 4'b0100; 
	if(x==?20'b??11?1?????1?0??111?) z |= 4'b0100; 
	if(x==?20'b?11?01?1????????111?) z |= 4'b0100; 
	if(x==?20'b?11??1?1???1?0???11?) z |= 4'b0100; 
	if(x==?20'b?11?111?1?????????11) z |= 4'b1000; 
	if(x==?20'b?1????10?????00?111?) z |= 4'b1000; 
	if(x==?20'b??????????1111??1?11) z |= 4'b0100; 
	if(x==?20'b?11?11??1????0??1?1?) z |= 4'b1000; 
	if(x==?20'b?11?11??1?????0?1?1?) z |= 4'b1000; 
	if(x==?20'b??1?01???????00?111?) z |= 4'b0100; 
	if(x==?20'b?????1???11??1?1?11?) z |= 4'b1000; 
	if(x==?20'b?1??11???10????0?1??) z |= 4'b1000; 
	if(x==?20'b??????1??11?1?1??11?) z |= 4'b0100; 
	if(x==?20'b?1??11???1?0???0?1??) z |= 4'b1000; 
	if(x==?20'b????????11????111?11) z |= 4'b1000; 
	if(x==?20'b?11???11???1?0??1?1?) z |= 4'b0100; 
	if(x==?20'b?11??111???1??????11) z |= 4'b0100; 
	if(x==?20'b?11??1??11???0??1??1) z |= 4'b1000; 
	if(x==?20'b??1???110?1?0????1??) z |= 4'b0100; 
	if(x==?20'b??1???11?01?0????1??) z |= 4'b0100; 
	if(x==?20'b?11???11???1??0?1?1?) z |= 4'b0100; 
	if(x==?20'b?11??1??11????0?1??1) z |= 4'b1000; 
	if(x==?20'b1???1?101????????1?1) z |= 4'b1000; 
	if(x==?20'b?1???111?????00?1??1) z |= 4'b0100; 
	if(x==?20'b1?1??????????1?1?111) z |= 4'b1000; 
	if(x==?20'b?1?1????????1?1??111) z |= 4'b0100; 
	if(x==?20'b???1?11?00??????1??1) z |= 4'b0100; 
	if(x==?20'b1????11???00????1??1) z |= 4'b1000; 
	if(x==?20'b??11??1??????00?1?11) z |= 4'b0100; 
	if(x==?20'b?11???1???11?0??1??1) z |= 4'b0100; 
	if(x==?20'b??11????????11??1?11) z |= 4'b0100; 
	if(x==?20'b?11???1???11??0?1??1) z |= 4'b0100; 
	if(x==?20'b????????11??11??1?1?) z |= 4'b0010; 
	if(x==?20'b????????1?1?1?1??11?) z |= 4'b0010; 
	if(x==?20'b???101?1???1?????1?1) z |= 4'b0100; 
	if(x==?20'b?11?1?1??1???0???11?) z |= 4'b1000; 
	if(x==?20'b?????????1?1?1?1?11?) z |= 4'b0001; 
	if(x==?20'b?1???11???11?0???11?) z |= 4'b0100; 
	if(x==?20'b????11????00?0??1??1) z |= 4'b1000; 
	if(x==?20'b????11????00??0?1??1) z |= 4'b1000; 
	if(x==?20'b??????1100???0??1??1) z |= 4'b0100; 
	if(x==?20'b??????1100????0?1??1) z |= 4'b0100; 
	if(x==?20'b?111?11??1??????11??) z |= 4'b0100; 
	if(x==?20'b111??11???1?????11??) z |= 4'b1000; 
	if(x==?20'b?11??1?1??1???0??11?) z |= 4'b0100; 
	if(x==?20'b?1??1??0?1?????0?1?1) z |= 4'b1000; 
	if(x==?20'b11????????????111?11) z |= 4'b1000; 
	if(x==?20'b??1?0??1??1?0????1?1) z |= 4'b0100; 
	if(x==?20'b111??11??????0???11?) z |= 4'b1000; 
	if(x==?20'b?111?11??????0???11?) z |= 4'b0100; 
	if(x==?20'b?11?111?1???????1?1?) z |= 4'b1000; 
	if(x==?20'b111??11???????0??11?) z |= 4'b1000; 
	if(x==?20'b?1??111?00??????1??1) z |= 4'b1100; 
	if(x==?20'b?111?11???????0??11?) z |= 4'b0100; 
	if(x==?20'b??1??111??00????1??1) z |= 4'b1100; 
	if(x==?20'b????11??????11??1??1) z |= 4'b0010; 
	if(x==?20'b11????1??????00?111?) z |= 4'b1000; 
	if(x==?20'b??11?1???????00?111?) z |= 4'b0100; 
	if(x==?20'b??????????11??111?1?) z |= 4'b0001; 
	if(x==?20'b??????11????11??1?11) z |= 4'b0100; 
	if(x==?20'b?11??111???1????1?1?) z |= 4'b0100; 
	if(x==?20'b?1???1?0?10???0??1??) z |= 4'b1000; 
	if(x==?20'b??1?0?1??01??0???1??) z |= 4'b0100; 
	if(x==?20'b?????????11?11??1?1?) z |= 4'b0010; 
	if(x==?20'b1?????1?1??1?1??11??) z |= 4'b1000; 
	if(x==?20'b???1?1??1??1?1??11??) z |= 4'b0100; 
	if(x==?20'b11??1??0?1???????1?1) z |= 4'b1000; 
	if(x==?20'b??????11??????111??1) z |= 4'b0001; 
	if(x==?20'b????11????????111?11) z |= 4'b1000; 
	if(x==?20'b1?1?111???0????????1) z |= 4'b1000; 
	if(x==?20'b??110??1??1??????1?1) z |= 4'b0100; 
	if(x==?20'b?????11?1?00????1??1) z |= 4'b1000; 
	if(x==?20'b1?????1?1??1??1?11??) z |= 4'b1000; 
	if(x==?20'b??1??10??10?????11??) z |= 4'b1000; 
	if(x==?20'b??1??01?01??????11??) z |= 4'b0100; 
	if(x==?20'b??1?1??1?1??1???11??) z |= 4'b0100; 
	if(x==?20'b?1??1??1?1??1???11??) z |= 4'b0100; 
	if(x==?20'b11??111????0???????1) z |= 4'b1000; 
	if(x==?20'b??11?1110??????????1) z |= 4'b0100; 
	if(x==?20'b???1?1??1??1??1?11??) z |= 4'b0100; 
	if(x==?20'b?1?1?111?0?????????1) z |= 4'b0100; 
	if(x==?20'b?11???1???????00111?) z |= 4'b1000; 
	if(x==?20'b?11??1??????00??111?) z |= 4'b0100; 
	if(x==?20'b?1??1??1??1?1???11??) z |= 4'b0100; 
	if(x==?20'b?11?111??1??????1?1?) z |= 4'b1000; 
	if(x==?20'b?1???01??01?????11??) z |= 4'b0100; 
	if(x==?20'b?????????11???111?1?) z |= 4'b0001; 
	if(x==?20'b?????11?00?1????1??1) z |= 4'b0100; 
	if(x==?20'b??11??1?0???0????11?) z |= 4'b0100; 
	if(x==?20'b????????11???11?1?11) z |= 4'b1000; 
	if(x==?20'b1???11???10?????11??) z |= 4'b1000; 
	if(x==?20'b11??1????1?????0?1?1) z |= 4'b1000; 
	if(x==?20'b?1???10???10????11??) z |= 4'b1000; 
	if(x==?20'b??1?1??1?1?????111??) z |= 4'b1000; 
	if(x==?20'b11???1?????0???0?11?) z |= 4'b1000; 
	if(x==?20'b??1?11????00????1??1) z |= 4'b1000; 
	if(x==?20'b?1??11????00????1??1) z |= 4'b1000; 
	if(x==?20'b??1???1??1??1?1??11?) z |= 4'b0100; 
	if(x==?20'b????1????100????111?) z |= 4'b1000; 
	if(x==?20'b?11??111??1?????1?1?) z |= 4'b0100; 
	if(x==?20'b1???11???1?0????11??) z |= 4'b1000; 
	if(x==?20'b??1?1??1??1????111??) z |= 4'b1000; 
	if(x==?20'b?1??1??1??1????111??) z |= 4'b1000; 
	if(x==?20'b?1?10???0????????111) z |= 4'b0100; 
	if(x==?20'b?1???1????1??1?1?11?) z |= 4'b1000; 
	if(x==?20'b??11???1??1?0????1?1) z |= 4'b0100; 
	if(x==?20'b???1??110?1?????11??) z |= 4'b0100; 
	if(x==?20'b??1??1??0??1?1???1?1) z |= 4'b0100; 
	if(x==?20'b???1??11?01?????11??) z |= 4'b0100; 
	if(x==?20'b1?1????0???0?????111) z |= 4'b1000; 
	if(x==?20'b??1??01?0????0???11?) z |= 4'b0100; 
	if(x==?20'b??????????11?11?1?11) z |= 4'b0100; 
	if(x==?20'b???????1001?????111?) z |= 4'b0100; 
	if(x==?20'b?1????1?1??0??1??1?1) z |= 4'b1000; 
	if(x==?20'b1???1???1??????011?1) z |= 4'b1000; 
	if(x==?20'b?1???10????0??0??11?) z |= 4'b1000; 
	if(x==?20'b1????1??1????0?0?1?1) z |= 4'b1000; 
	if(x==?20'b??1?1?1?1?1??1???1??) z |= 4'b0100; 
	if(x==?20'b??1?1?1??1?1?1???1??) z |= 4'b0100; 
	if(x==?20'b??1??1?11?1??1???1??) z |= 4'b0100; 
	if(x==?20'b?1????1?1????00?111?) z |= 4'b1000; 
	if(x==?20'b???1???1???10???11?1) z |= 4'b0100; 
	if(x==?20'b???1??1????10?0??1?1) z |= 4'b0100; 
	if(x==?20'b??1??1?1?1?1?1???1??) z |= 4'b0100; 
	if(x==?20'b???1???110??????111?) z |= 4'b0100; 
	if(x==?20'b?1??1?1?1?1???1??1??) z |= 4'b1000; 
	if(x==?20'b1???1?????01????111?) z |= 4'b1000; 
	if(x==?20'b1???111???0???????11) z |= 4'b1000; 
	if(x==?20'b??1???11?0??0???1??1) z |= 4'b0100; 
	if(x==?20'b11???????????11?1?11) z |= 4'b1000; 
	if(x==?20'b?1??1?1??1?1??1??1??) z |= 4'b1000; 
	if(x==?20'b??11?????????11?1?11) z |= 4'b0100; 
	if(x==?20'b??1??1?????1?00?111?) z |= 4'b0100; 
	if(x==?20'b?1???1?11?1???1??1??) z |= 4'b1000; 
	if(x==?20'b????????11???11?1?1?) z |= 4'b0010; 
	if(x==?20'b1??????011???????111) z |= 4'b1000; 
	if(x==?20'b?1???1?1?1?1??1??1??) z |= 4'b1000; 
	if(x==?20'b1?1??1?????1???111??) z |= 4'b1000; 
	if(x==?20'b???1?111?0????????11) z |= 4'b0100; 
	if(x==?20'b?1??11?0???????01??1) z |= 4'b1000; 
	if(x==?20'b??1?0?11????0???1??1) z |= 4'b0100; 
	if(x==?20'b?1??1??011???????1?1) z |= 4'b1000; 
	if(x==?20'b??????????11?11?1?1?) z |= 4'b0001; 
	if(x==?20'b???10?????11?????111) z |= 4'b0100; 
	if(x==?20'b???1?111?0??????1??1) z |= 4'b0100; 
	if(x==?20'b??1?111?1?0????????1) z |= 4'b1000; 
	if(x==?20'b??1???110???0????11?) z |= 4'b0100; 
	if(x==?20'b?1??111?1??0???????1) z |= 4'b1000; 
	if(x==?20'b?1??11?????0???0?11?) z |= 4'b1000; 
	if(x==?20'b1?1?1?10?????????1?1) z |= 4'b1000; 
	if(x==?20'b????0?11?0??????1?11) z |= 4'b0100; 
	if(x==?20'b????1?1?1?1??1???1??) z |= 4'b0010; 
	if(x==?20'b??1?1?1??11??1???1??) z |= 4'b0100; 
	if(x==?20'b??1?0??1??11?????1?1) z |= 4'b0100; 
	if(x==?20'b?1?101?1?????????1?1) z |= 4'b0100; 
	if(x==?20'b?1??1???11?????0?1?1) z |= 4'b1000; 
	if(x==?20'b????11???????11?1??1) z |= 4'b0010; 
	if(x==?20'b??1??1110??1???????1) z |= 4'b0100; 
	if(x==?20'b??1??1?1?11??1???1??) z |= 4'b0100; 
	if(x==?20'b?1???111?0?1???????1) z |= 4'b0100; 
	if(x==?20'b??????11?????11?1??1) z |= 4'b0001; 
	if(x==?20'b?1???1??1??0???0?11?) z |= 4'b1000; 
	if(x==?20'b????11???????11?1?11) z |= 4'b1000; 
	if(x==?20'b??11??11?0??????1??1) z |= 4'b0100; 
	if(x==?20'b??1???1?0??10????11?) z |= 4'b0100; 
	if(x==?20'b??????11?????11?1?11) z |= 4'b0100; 
	if(x==?20'b?1??1?1??11???1??1??) z |= 4'b1000; 
	if(x==?20'b?1???1?1?11???1??1??) z |= 4'b1000; 
	if(x==?20'b11??11?0????????1??1) z |= 4'b1000; 
	if(x==?20'b??110?11????????1??1) z |= 4'b0100; 
	if(x==?20'b?1??11???10??0???1??) z |= 4'b1000; 
	if(x==?20'b?????1?1?1?1??1??1??) z |= 4'b0001; 
	if(x==?20'b??1????1??110????1?1) z |= 4'b0100; 
	if(x==?20'b?????110?????0?0?1?1) z |= 4'b1000; 
	if(x==?20'b????011?????0?0??1?1) z |= 4'b0100; 
	if(x==?20'b?1???1111?0?????1??1) z |= 4'b1100; 
	if(x==?20'b1???1????????0?011?1) z |= 4'b1000; 
	if(x==?20'b?1??11???1?0?0???1??) z |= 4'b1000; 
	if(x==?20'b?1??11???1?0??0??1??) z |= 4'b1000; 
	if(x==?20'b???1??1?????000??1?1) z |= 4'b0100; 
	if(x==?20'b??1???110?1??0???1??) z |= 4'b0100; 
	if(x==?20'b1?1??1??1??????0?1?1) z |= 4'b1000; 
	if(x==?20'b???1???1????0?0?11?1) z |= 4'b0100; 
	if(x==?20'b1????1???????000?1?1) z |= 4'b1000; 
	if(x==?20'b??1???110?1???0??1??) z |= 4'b0100; 
	if(x==?20'b??1???11?01???0??1??) z |= 4'b0100; 
	if(x==?20'b?1??1?1????1???111??) z |= 4'b1000; 
	if(x==?20'b??11??110????????11?) z |= 4'b0100; 
	if(x==?20'b??1??1??1??11???11??) z |= 4'b0100; 
	if(x==?20'b?1???1??1??11???11??) z |= 4'b0100; 
	if(x==?20'b1???????1?????0011?1) z |= 4'b1000; 
	if(x==?20'b?1?1??1????10????1?1) z |= 4'b0100; 
	if(x==?20'b11??11?????0?????11?) z |= 4'b1000; 
	if(x==?20'b11??11?????????01??1) z |= 4'b1000; 
	if(x==?20'b?11???1?1?????0?111?) z |= 4'b1000; 
	if(x==?20'b?????????11??11?1?1?) z |= 4'b0011; 
	if(x==?20'b??11??11????0???1??1) z |= 4'b0100; 
	if(x==?20'b????111?1?0???????11) z |= 4'b1000; 
	if(x==?20'b???1???????100??11?1) z |= 4'b0100; 
	if(x==?20'b11??1???11???????1?1) z |= 4'b1000; 
	if(x==?20'b??1???1?1??1???111??) z |= 4'b1000; 
	if(x==?20'b?1????1?1??1???111??) z |= 4'b1000; 
	if(x==?20'b11???1??1??0?????11?) z |= 4'b1000; 
	if(x==?20'b?11??1?????1?0??111?) z |= 4'b0100; 
	if(x==?20'b??????11011??????11?) z |= 4'b0100; 
	if(x==?20'b????11???110?????11?) z |= 4'b1000; 
	if(x==?20'b??11??1?0??1?????11?) z |= 4'b0100; 
	if(x==?20'b1?1???10?1???????1?1) z |= 4'b1000; 
	if(x==?20'b?????111?0?1??????11) z |= 4'b0100; 
	if(x==?20'b?1?1?1????1??1???1?1) z |= 4'b0100; 
	if(x==?20'b????1?1??1???0?0?1?1) z |= 4'b1000; 
	if(x==?20'b??1???1???1?01???11?) z |= 4'b0100; 
	if(x==?20'b?1?1??1?1????1??11??) z |= 4'b0100; 
	if(x==?20'b???1??11?0??????1?11) z |= 4'b0100; 
	if(x==?20'b??1?0?1?0????0???11?) z |= 4'b0100; 
	if(x==?20'b?1?101????1??????1?1) z |= 4'b0100; 
	if(x==?20'b1?1???1??1????1??1?1) z |= 4'b1000; 
	if(x==?20'b??11???1??11?????1?1) z |= 4'b0100; 
	if(x==?20'b?1??1??0?1???0???1?1) z |= 4'b1000; 
	if(x==?20'b11??11?????????0?11?) z |= 4'b1000; 
	if(x==?20'b?1???1?0???0??0??11?) z |= 4'b1000; 
	if(x==?20'b1???11??11???????11?) z |= 4'b1000; 
	if(x==?20'b?????111?0?1????1??1) z |= 4'b0100; 
	if(x==?20'b??11??11????0????11?) z |= 4'b0100; 
	if(x==?20'b1???11?0????????1?11) z |= 4'b1000; 
	if(x==?20'b?1???1???1????10?11?) z |= 4'b1000; 
	if(x==?20'b?????1?1??1?0?0??1?1) z |= 4'b0100; 
	if(x==?20'b???10?11????????1?11) z |= 4'b0100; 
	if(x==?20'b??1?1?101????????1?1) z |= 4'b1000; 
	if(x==?20'b?11?0110????????1??1) z |= 4'b1100; 
	if(x==?20'b1???11??1?1??????11?) z |= 4'b1000; 
	if(x==?20'b?1?1??1?1?????1?11??) z |= 4'b0100; 
	if(x==?20'b??1?0??1??1???0??1?1) z |= 4'b0100; 
	if(x==?20'b1?1?1??0?????????111) z |= 4'b1000; 
	if(x==?20'b11???1??1??????0?11?) z |= 4'b1000; 
	if(x==?20'b1?1?????1??0?????111) z |= 4'b1000; 
	if(x==?20'b?1?10??1?????????111) z |= 4'b0100; 
	if(x==?20'b???1?01??????0??111?) z |= 4'b0100; 
	if(x==?20'b???1??11?1?1?????11?) z |= 4'b0100; 
	if(x==?20'b??1??11?00??????1??1) z |= 4'b0100; 
	if(x==?20'b?1???11???00????1??1) z |= 4'b1000; 
	if(x==?20'b?11???1??????00?1?11) z |= 4'b0100; 
	if(x==?20'b?11??1???????00?1?11) z |= 4'b1000; 
	if(x==?20'b?????111111????????1) z |= 4'b0100; 
	if(x==?20'b1????10???????0?111?) z |= 4'b1000; 
	if(x==?20'b1?1??1?????1??1?11??) z |= 4'b1000; 
	if(x==?20'b?1?1????0??1?????111) z |= 4'b0100; 
	if(x==?20'b?11?????????11??1?11) z |= 4'b0100; 
	if(x==?20'b??11??1????10????11?) z |= 4'b0100; 
	if(x==?20'b???1??11??11?????11?) z |= 4'b0100; 
	if(x==?20'b11?????01????????111) z |= 4'b1000; 
	if(x==?20'b?1??1????1???0?0?1?1) z |= 4'b1000; 
	if(x==?20'b?1??01?1???1?????1?1) z |= 4'b0100; 
	if(x==?20'b????111??111???????1) z |= 4'b1000; 
	if(x==?20'b?1??1110?1???????1??) z |= 4'b1000; 
	if(x==?20'b?1??11?01???????1??1) z |= 4'b1000; 
	if(x==?20'b??1???11?0?1????1??1) z |= 4'b0100; 
	if(x==?20'b??1??111??1??1???1??) z |= 4'b0100; 
	if(x==?20'b??110??????1?????111) z |= 4'b0100; 
	if(x==?20'b??1????1??1?0?0??1?1) z |= 4'b0100; 
	if(x==?20'b????11???????000?1?1) z |= 4'b1000; 
	if(x==?20'b?1?1??1??1???1???11?) z |= 4'b0100; 
	if(x==?20'b??????11????000??1?1) z |= 4'b0100; 
	if(x==?20'b??1?0111??1??????1??) z |= 4'b0100; 
	if(x==?20'b????1???1????0?011?1) z |= 4'b1000; 
	if(x==?20'b??1??11?1?1??1???1??) z |= 4'b0100; 
	if(x==?20'b1?1??1???10?????11??) z |= 4'b1000; 
	if(x==?20'b??11??1???1??1???11?) z |= 4'b0100; 
	if(x==?20'b??1?0?11???1????1??1) z |= 4'b0100; 
	if(x==?20'b??1??11??1?1?1???1??) z |= 4'b0100; 
	if(x==?20'b?????1??1????000?1?1) z |= 4'b1000; 
	if(x==?20'b1?1?1??????????011?1) z |= 4'b1000; 
	if(x==?20'b1?1??1???1?0????11??) z |= 4'b1000; 
	if(x==?20'b?11???????????111?11) z |= 4'b1000; 
	if(x==?20'b?1?1??1?0?1?????11??) z |= 4'b0100; 
	if(x==?20'b?1?1??1??01?????11??) z |= 4'b0100; 
	if(x==?20'b11???1???1????1??11?) z |= 4'b1000; 
	if(x==?20'b?1?1???1????0???11?1) z |= 4'b0100; 
	if(x==?20'b?1?1??1?????0?0??1?1) z |= 4'b0100; 
	if(x==?20'b1?1??1???????0?0?1?1) z |= 4'b1000; 
	if(x==?20'b?1??11??1??0?????11?) z |= 4'b1000; 
	if(x==?20'b?1??11??1??????01??1) z |= 4'b1000; 
	if(x==?20'b?1???11?1?1???1??1??) z |= 4'b1000; 
	if(x==?20'b??????1????1000??1?1) z |= 4'b0100; 
	if(x==?20'b???????1???10?0?11?1) z |= 4'b0100; 
	if(x==?20'b??1?????0???0?0??111) z |= 4'b0100; 
	if(x==?20'b1?1??1????1???1??11?) z |= 4'b1000; 
	if(x==?20'b?1???11??1?1??1??1??) z |= 4'b1000; 
	if(x==?20'b?1?????????0?0?0?111) z |= 4'b1000; 
	if(x==?20'b11??????1??????011?1) z |= 4'b1000; 
	if(x==?20'b??1???110??1?????11?) z |= 4'b0100; 
	if(x==?20'b?11???1??????00?111?) z |= 4'b1000; 
	if(x==?20'b?1??11?????1???01??1) z |= 4'b1000; 
	if(x==?20'b?11??1???????00?111?) z |= 4'b0100; 
	if(x==?20'b????111???0???0???11) z |= 4'b1000; 
	if(x==?20'b??1???11???10???1??1) z |= 4'b0100; 
	if(x==?20'b??11??1?0????0???11?) z |= 4'b0100; 
	if(x==?20'b??11??1?0?????0??11?) z |= 4'b0100; 
	if(x==?20'b11??1????1???0???1?1) z |= 4'b1000; 
	if(x==?20'b??11???????10???11?1) z |= 4'b0100; 
	if(x==?20'b1?1?1????1????0??1?1) z |= 4'b1000; 
	if(x==?20'b1???111?1???????1??1) z |= 4'b1000; 
	if(x==?20'b?????111?0???0????11) z |= 4'b0100; 
	if(x==?20'b11???1?????0?0???11?) z |= 4'b1000; 
	if(x==?20'b??1??1?11????1??11??) z |= 4'b0100; 
	if(x==?20'b1???11?????????0111?) z |= 4'b1000; 
	if(x==?20'b11???1?????0??0??11?) z |= 4'b1000; 
	if(x==?20'b???1??11????0???111?) z |= 4'b0100; 
	if(x==?20'b1?1?1?1?1????????1?1) z |= 4'b1000; 
	if(x==?20'b?1?1???1??1??0???1?1) z |= 4'b0100; 
	if(x==?20'b??1???110?1?????1??1) z |= 4'b0100; 
	if(x==?20'b?1????110?1?????1??1) z |= 4'b0100; 
	if(x==?20'b??11???1??1???0??1?1) z |= 4'b0100; 
	if(x==?20'b????1????1???0?0?111) z |= 4'b1000; 
	if(x==?20'b1???111????1????1??1) z |= 4'b1000; 
	if(x==?20'b?1??11?0?1??????1??1) z |= 4'b1000; 
	if(x==?20'b1????1??1??????0111?) z |= 4'b1000; 
	if(x==?20'b?1??11??1??????0?11?) z |= 4'b1000; 
	if(x==?20'b1???1???1????0??11?1) z |= 4'b1000; 
	if(x==?20'b???1?111???1????1??1) z |= 4'b0100; 
	if(x==?20'b??1???1?1??1?1??11??) z |= 4'b1000; 
	if(x==?20'b??1??1?11?????1?11??) z |= 4'b0100; 
	if(x==?20'b????11?01???????1?11) z |= 4'b1000; 
	if(x==?20'b??????11?0?1????1?11) z |= 4'b0100; 
	if(x==?20'b?1???1??1??1?1??11??) z |= 4'b0100; 
	if(x==?20'b?11?1??0?1???????1?1) z |= 4'b1000; 
	if(x==?20'b?1??1?1????1??1?11??) z |= 4'b1000; 
	if(x==?20'b??1?0?11??1?????1??1) z |= 4'b0100; 
	if(x==?20'b???????1??1?0?0??111) z |= 4'b0100; 
	if(x==?20'b???1??1????10???111?) z |= 4'b0100; 
	if(x==?20'b?1?1?1?1???1?????1?1) z |= 4'b0100; 
	if(x==?20'b??1???11???10????11?) z |= 4'b0100; 
	if(x==?20'b????11?0???1????1?11) z |= 4'b1000; 
	if(x==?20'b?1??11??1??????011??) z |= 4'b1000; 
	if(x==?20'b11??111??1???????1??) z |= 4'b1000; 
	if(x==?20'b?11?0??1??1??????1?1) z |= 4'b0100; 
	if(x==?20'b11??11??1???????1??1) z |= 4'b1000; 
	if(x==?20'b????0?11???1????1?11) z |= 4'b0100; 
	if(x==?20'b??11?11??0??????1??1) z |= 4'b0100; 
	if(x==?20'b??1???1?1??1??1?11??) z |= 4'b1000; 
	if(x==?20'b?1????1?1??1??1?11??) z |= 4'b1000; 
	if(x==?20'b???1???1???1??0?11?1) z |= 4'b0100; 
	if(x==?20'b?11?111????0???????1) z |= 4'b1000; 
	if(x==?20'b?11??1110??????????1) z |= 4'b0100; 
	if(x==?20'b?1???1??1??1??1?11??) z |= 4'b0100; 
	if(x==?20'b??11?111??1??????1??) z |= 4'b0100; 
	if(x==?20'b??1???11???10???11??) z |= 4'b0100; 
	if(x==?20'b11??11?????1????1??1) z |= 4'b1000; 
	if(x==?20'b??1???11?0???0??1??1) z |= 4'b0100; 
	if(x==?20'b?11???1?0???0????11?) z |= 4'b0100; 
	if(x==?20'b111??1????0???????11) z |= 4'b1000; 
	if(x==?20'b11???110????????1??1) z |= 4'b1000; 
	if(x==?20'b??11011?????????1??1) z |= 4'b0100; 
	if(x==?20'b??1???11?0????0?1??1) z |= 4'b0100; 
	if(x==?20'b??11??11???1????1??1) z |= 4'b0100; 
	if(x==?20'b?11?1????1?????0?1?1) z |= 4'b1000; 
	if(x==?20'b?111??1??0????????11) z |= 4'b0100; 
	if(x==?20'b?11??1?????0???0?11?) z |= 4'b1000; 
	if(x==?20'b??1?11???1?0????11??) z |= 4'b1000; 
	if(x==?20'b?1??11?0?????0??1??1) z |= 4'b1000; 
	if(x==?20'b?1??11?0??????0?1??1) z |= 4'b1000; 
	if(x==?20'b?????10?1?????0?111?) z |= 4'b1010; 
	if(x==?20'b?1??1?1??????0?0?1?1) z |= 4'b1000; 
	if(x==?20'b??1?0?11?????0??1??1) z |= 4'b0100; 
	if(x==?20'b?11????1??1?0????1?1) z |= 4'b0100; 
	if(x==?20'b??1?0?11??????0?1??1) z |= 4'b0100; 
	if(x==?20'b?1????110?1?????11??) z |= 4'b0100; 
	if(x==?20'b?????01????1?0??111?) z |= 4'b0101; 
	if(x==?20'b??1??1?1????0?0??1?1) z |= 4'b0100; 
	if(x==?20'b??1?1???1??????011?1) z |= 4'b1000; 
	if(x==?20'b11??11??1????????11?) z |= 4'b1000; 
	if(x==?20'b??1???1???11?1???11?) z |= 4'b0100; 
	if(x==?20'b?1???1??11????1??11?) z |= 4'b1000; 
	if(x==?20'b??1??1??1????0?0?1?1) z |= 4'b1000; 
	if(x==?20'b1?1???1?11???????1?1) z |= 4'b1000; 
	if(x==?20'b??1???110?????0??11?) z |= 4'b0100; 
	if(x==?20'b?1??11?????0?0???11?) z |= 4'b1000; 
	if(x==?20'b??11??11???1?????11?) z |= 4'b0100; 
	if(x==?20'b?????1??11?0????1?11) z |= 4'b1000; 
	if(x==?20'b?1?????1???10???11?1) z |= 4'b0100; 
	if(x==?20'b?1????1????10?0??1?1) z |= 4'b0100; 
	if(x==?20'b?1??11????????001??1) z |= 4'b1000; 
	if(x==?20'b??1???11????00??1??1) z |= 4'b0100; 
	if(x==?20'b???10?1??????0??111?) z |= 4'b0100; 
	if(x==?20'b?1?????110??????111?) z |= 4'b0100; 
	if(x==?20'b?1??1???11???0???1?1) z |= 4'b1000; 
	if(x==?20'b1????1?0??????0?111?) z |= 4'b1000; 
	if(x==?20'b??1?1?????01????111?) z |= 4'b1000; 
	if(x==?20'b?1???1??1??0?0???11?) z |= 4'b1000; 
	if(x==?20'b??1?111???0???????11) z |= 4'b1000; 
	if(x==?20'b??????1?0?11????1?11) z |= 4'b0100; 
	if(x==?20'b??1??110?1???0???11?) z |= 4'b1100; 
	if(x==?20'b????11??1??????0111?) z |= 4'b1000; 
	if(x==?20'b?1???1??1??0??0??11?) z |= 4'b1000; 
	if(x==?20'b??1????11????1??111?) z |= 4'b0100; 
	if(x==?20'b1???111??1???????11?) z |= 4'b1000; 
	if(x==?20'b?111??1?0????????11?) z |= 4'b0100; 
	if(x==?20'b1???11??1???????1?11) z |= 4'b1000; 
	if(x==?20'b??1???1?0??1?0???11?) z |= 4'b0100; 
	if(x==?20'b111?1????1???????1?1) z |= 4'b1000; 
	if(x==?20'b??1???1?0??1??0??11?) z |= 4'b0100; 
	if(x==?20'b?1?1?1????11?????1?1) z |= 4'b0100; 
	if(x==?20'b?1??111????0??????11) z |= 4'b1000; 
	if(x==?20'b?1??011???1???0??11?) z |= 4'b1100; 
	if(x==?20'b??1??1110?????????11) z |= 4'b0100; 
	if(x==?20'b?1???111?0????????11) z |= 4'b0100; 
	if(x==?20'b111??1?????0?????11?) z |= 4'b1000; 
	if(x==?20'b1?1?1???1????????111) z |= 4'b1000; 
	if(x==?20'b????111?1??1????1??1) z |= 4'b1000; 
	if(x==?20'b???1?111??1??????11?) z |= 4'b0100; 
	if(x==?20'b1???11?????1????1?11) z |= 4'b1000; 
	if(x==?20'b??????11???10???111?) z |= 4'b0100; 
	if(x==?20'b?111???1??1??????1?1) z |= 4'b0100; 
	if(x==?20'b???1??11???1????1?11) z |= 4'b0100; 
	if(x==?20'b??1????1??11??0??1?1) z |= 4'b0100; 
	if(x==?20'b1?1?1???1???????11?1) z |= 4'b1000; 
	if(x==?20'b?1??1??????1??1?111?) z |= 4'b1000; 
	if(x==?20'b?1?1???1???1?????111) z |= 4'b0100; 
	if(x==?20'b1?1??1??1????0???1?1) z |= 4'b1000; 
	if(x==?20'b?1??111?11???????1??) z |= 4'b1000; 
	if(x==?20'b11???1????0?????1?11) z |= 4'b1000; 
	if(x==?20'b?1?11?1??1???????11?) z |= 4'b0100; 
	if(x==?20'b??11??1??0??????1?11) z |= 4'b0100; 
	if(x==?20'b1?1?11???1???????11?) z |= 4'b1000; 
	if(x==?20'b?1????1??1???0?0?1?1) z |= 4'b1000; 
	if(x==?20'b?1?1??11?1???????11?) z |= 4'b0100; 
	if(x==?20'b1???????1????00?11?1) z |= 4'b1000; 
	if(x==?20'b1?1?1?1???1??????11?) z |= 4'b1000; 
	if(x==?20'b?1?1?1?1?1???????11?) z |= 4'b0100; 
	if(x==?20'b11??11???????0??1??1) z |= 4'b1000; 
	if(x==?20'b1?1?11????1??????11?) z |= 4'b1000; 
	if(x==?20'b?1?1???1???1????11?1) z |= 4'b0100; 
	if(x==?20'b?1?1??1????1??0??1?1) z |= 4'b0100; 
	if(x==?20'b11??11????????0?1??1) z |= 4'b1000; 
	if(x==?20'b?1??11??1??1????1??1) z |= 4'b1000; 
	if(x==?20'b??11??11?????0??1??1) z |= 4'b0100; 
	if(x==?20'b?1?1??11??1??????11?) z |= 4'b0100; 
	if(x==?20'b?1???1101???????1??1) z |= 4'b1000; 
	if(x==?20'b??11??11??????0?1??1) z |= 4'b0100; 
	if(x==?20'b1?1??1?1??1??????11?) z |= 4'b1000; 
	if(x==?20'b??1??1????1?0?0??1?1) z |= 4'b0100; 
	if(x==?20'b??110?1?????????1?11) z |= 4'b0100; 
	if(x==?20'b11???1?0????????1?11) z |= 4'b1000; 
	if(x==?20'b???1???????1?00?11?1) z |= 4'b0100; 
	if(x==?20'b??11??11?1??????11??) z |= 4'b0100; 
	if(x==?20'b??1??111??11?????1??) z |= 4'b0100; 
	if(x==?20'b?11???11?0??????1??1) z |= 4'b0100; 
	if(x==?20'b1???11??1???????111?) z |= 4'b1000; 
	if(x==?20'b11??11????1?????11??) z |= 4'b1000; 
	if(x==?20'b111????0?????????111) z |= 4'b1000; 
	if(x==?20'b?1???110???1????1??1) z |= 4'b1000; 
	if(x==?20'b?1110????????????111) z |= 4'b0100; 
	if(x==?20'b??1?011????1????1??1) z |= 4'b0100; 
	if(x==?20'b?1??111????0?????11?) z |= 4'b1000; 
	if(x==?20'b??1??1110????????11?) z |= 4'b0100; 
	if(x==?20'b?1??1????????0?0?111) z |= 4'b1000; 
	if(x==?20'b?11?11?0????????1??1) z |= 4'b1000; 
	if(x==?20'b?11?0?11????????1??1) z |= 4'b0100; 
	if(x==?20'b??1????1????0?0??111) z |= 4'b0100; 
	if(x==?20'b11???1??1?1?????11??) z |= 4'b1000; 
	if(x==?20'b???1??11???1????111?) z |= 4'b0100; 
	if(x==?20'b??1???1???1??10??11?) z |= 4'b0100; 
	if(x==?20'b??11??1??1?1????11??) z |= 4'b0100; 
	if(x==?20'b??1?1????????0?011?1) z |= 4'b1000; 
	if(x==?20'b11??11???????0???11?) z |= 4'b1000; 
	if(x==?20'b11??11????????0??11?) z |= 4'b1000; 
	if(x==?20'b??11??11?????0???11?) z |= 4'b0100; 
	if(x==?20'b?1???1???1???01??11?) z |= 4'b1000; 
	if(x==?20'b?1????1?????000??1?1) z |= 4'b0100; 
	if(x==?20'b??11??11??????0??11?) z |= 4'b0100; 
	if(x==?20'b?1?????1????0?0?11?1) z |= 4'b0100; 
	if(x==?20'b??1??1???????000?1?1) z |= 4'b1000; 
	if(x==?20'b11??1???1???????111?) z |= 4'b1000; 
	if(x==?20'b?1??111??1????0????1) z |= 4'b1000; 
	if(x==?20'b?1??????1????0?011?1) z |= 4'b1000; 
	if(x==?20'b11???1??1????0???11?) z |= 4'b1000; 
	if(x==?20'b?11???110????????11?) z |= 4'b0100; 
	if(x==?20'b??1?????1?????0011?1) z |= 4'b1000; 
	if(x==?20'b11???1??1?????0??11?) z |= 4'b1000; 
	if(x==?20'b?11?11?????0?????11?) z |= 4'b1000; 
	if(x==?20'b?11?11?????????01??1) z |= 4'b1000; 
	if(x==?20'b?????1?01?????0?111?) z |= 4'b1000; 
	if(x==?20'b?1??1?????0???0?111?) z |= 4'b1000; 
	if(x==?20'b?11???11????0???1??1) z |= 4'b0100; 
	if(x==?20'b??1??111??1??0?????1) z |= 4'b0100; 
	if(x==?20'b????111?11???????11?) z |= 4'b1000; 
	if(x==?20'b??1????1?0???0??111?) z |= 4'b0100; 
	if(x==?20'b??11??1????1?0???11?) z |= 4'b0100; 
	if(x==?20'b????0?1????1?0??111?) z |= 4'b0100; 
	if(x==?20'b?11?1???11???????1?1) z |= 4'b1000; 
	if(x==?20'b?1?????????100??11?1) z |= 4'b0100; 
	if(x==?20'b??11???1???1????111?) z |= 4'b0100; 
	if(x==?20'b??11??1????1??0??11?) z |= 4'b0100; 
	if(x==?20'b??1????????10?0?11?1) z |= 4'b0100; 
	if(x==?20'b?11??1??1??0?????11?) z |= 4'b1000; 
	if(x==?20'b??11????11??????1?11) z |= 4'b0100; 
	if(x==?20'b????11??1??1????1?11) z |= 4'b1000; 
	if(x==?20'b?11???1?0??1?????11?) z |= 4'b0100; 
	if(x==?20'b1?1?111?????????1??1) z |= 4'b1000; 
	if(x==?20'b??1?011???1?????1??1) z |= 4'b0100; 
	if(x==?20'b?1?1?111????????1??1) z |= 4'b0100; 
	if(x==?20'b?????111??11?????11?) z |= 4'b0100; 
	if(x==?20'b?1????11?0??????1?11) z |= 4'b0100; 
	if(x==?20'b?11????1??11?????1?1) z |= 4'b0100; 
	if(x==?20'b11???11?1???????1??1) z |= 4'b1000; 
	if(x==?20'b?1?1??1?????0???111?) z |= 4'b0100; 
	if(x==?20'b11????????11????1?11) z |= 4'b1000; 
	if(x==?20'b1?1??1?????????0111?) z |= 4'b1000; 
	if(x==?20'b?11?11?????????0?11?) z |= 4'b1000; 
	if(x==?20'b1?1?1????????0??11?1) z |= 4'b1000; 
	if(x==?20'b??1?11??11???????11?) z |= 4'b1000; 
	if(x==?20'b?11???11????0????11?) z |= 4'b0100; 
	if(x==?20'b??1?11?0????????1?11) z |= 4'b1000; 
	if(x==?20'b?1??0?11????????1?11) z |= 4'b0100; 
	if(x==?20'b?1??11??1????0??1??1) z |= 4'b1000; 
	if(x==?20'b??1?11??1?1??????11?) z |= 4'b1000; 
	if(x==?20'b?1?1???1??????0?11?1) z |= 4'b0100; 
	if(x==?20'b????????????111???11) z |= 4'b0010; 
	if(x==?20'b?1??11??1?????0?1??1) z |= 4'b1000; 
	if(x==?20'b11???11????1????1??1) z |= 4'b1000; 
	if(x==?20'b??11?11????1????1??1) z |= 4'b0100; 
	if(x==?20'b?11??1??1??????0?11?) z |= 4'b1000; 
	if(x==?20'b11??????1????0??11?1) z |= 4'b1000; 
	if(x==?20'b?1???110?1???????11?) z |= 4'b1000; 
	if(x==?20'b1?1?????1?????0?11?1) z |= 4'b1000; 
	if(x==?20'b?1???01??????0??111?) z |= 4'b0100; 
	if(x==?20'b?1????11?1?1?????11?) z |= 4'b0100; 
	if(x==?20'b111?11??????????1??1) z |= 4'b1000; 
	if(x==?20'b?1??11?????1?0??1??1) z |= 4'b1000; 
	if(x==?20'b??1??10???????0?111?) z |= 4'b1000; 
	if(x==?20'b?111??11????????1??1) z |= 4'b0100; 
	if(x==?20'b?1??11?????1??0?1??1) z |= 4'b1000; 
	if(x==?20'b11??111??????????11?) z |= 4'b1000; 
	if(x==?20'b??1?011???1??????11?) z |= 4'b0100; 
	if(x==?20'b??1???11???1?0??1??1) z |= 4'b0100; 
	if(x==?20'b?11???1????10????11?) z |= 4'b0100; 
	if(x==?20'b?1????11??11?????11?) z |= 4'b0100; 
	if(x==?20'b?????????????111??11) z |= 4'b0001; 
	if(x==?20'b??1???11???1??0?1??1) z |= 4'b0100; 
	if(x==?20'b??11?111?????????11?) z |= 4'b0100; 
	if(x==?20'b?1?1???????1?0??11?1) z |= 4'b0100; 
	if(x==?20'b??11???????1??0?11?1) z |= 4'b0100; 
	if(x==?20'b1???11???????0??111?) z |= 4'b1000; 
	if(x==?20'b??????1111??????1?11) z |= 4'b1000; 
	if(x==?20'b???1??11??????0?111?) z |= 4'b0100; 
	if(x==?20'b1????1??1????0??111?) z |= 4'b1000; 
	if(x==?20'b?1??11??1????0???11?) z |= 4'b1000; 
	if(x==?20'b1????1??1?????0?111?) z |= 4'b1000; 
	if(x==?20'b?11???1???1??1???11?) z |= 4'b0100; 
	if(x==?20'b????11????11????1?11) z |= 4'b0100; 
	if(x==?20'b???1??1????1?0??111?) z |= 4'b0100; 
	if(x==?20'b111?11???????????11?) z |= 4'b1000; 
	if(x==?20'b???1??1????1??0?111?) z |= 4'b0100; 
	if(x==?20'b?111??11?????????11?) z |= 4'b0100; 
	if(x==?20'b?11??1???1????1??11?) z |= 4'b1000; 
	if(x==?20'b?1??11??1????0??11??) z |= 4'b1000; 
	if(x==?20'b??1???11???1??0??11?) z |= 4'b0100; 
	if(x==?20'b?11?????1??????011?1) z |= 4'b1000; 
	if(x==?20'b111??1??1????????11?) z |= 4'b1000; 
	if(x==?20'b????1?1??????1?1?1?1) z |= 4'b1000; 
	if(x==?20'b??1???11???1??0?11??) z |= 4'b0100; 
	if(x==?20'b?11???1?0?????0??11?) z |= 4'b0100; 
	if(x==?20'b?111??1????1?????11?) z |= 4'b0100; 
	if(x==?20'b?11?1????1???0???1?1) z |= 4'b1000; 
	if(x==?20'b?11????????10???11?1) z |= 4'b0100; 
	if(x==?20'b??1?111?1???????1??1) z |= 4'b1000; 
	if(x==?20'b?11??1?????0?0???11?) z |= 4'b1000; 
	if(x==?20'b??1?11?????????0111?) z |= 4'b1000; 
	if(x==?20'b?????1?1????1?1??1?1) z |= 4'b0100; 
	if(x==?20'b1?1?11??????????1?11) z |= 4'b1000; 
	if(x==?20'b?1????11????0???111?) z |= 4'b0100; 
	if(x==?20'b??1111??????????1?11) z |= 4'b0100; 
	if(x==?20'b????11??11??????1?1?) z |= 4'b0010; 
	if(x==?20'b11????11????????1?11) z |= 4'b1000; 
	if(x==?20'b?1?1??11????????1?11) z |= 4'b0100; 
	if(x==?20'b?11????1??1???0??1?1) z |= 4'b0100; 
	if(x==?20'b??1?111????1????1??1) z |= 4'b1000; 
	if(x==?20'b??1??1??1??????0111?) z |= 4'b1000; 
	if(x==?20'b??1?1???1????0??11?1) z |= 4'b1000; 
	if(x==?20'b?1???111???1????1??1) z |= 4'b0100; 
	if(x==?20'b?1?1?11??1???????11?) z |= 4'b0100; 
	if(x==?20'b11???1??1???????1?11) z |= 4'b1000; 
	if(x==?20'b????111???00???????1) z |= 4'b1000; 
	if(x==?20'b????1?1?????1?1??1?1) z |= 4'b0110; 
	if(x==?20'b??1??110?????0??111?) z |= 4'b1100; 
	if(x==?20'b?????11100?????????1) z |= 4'b0100; 
	if(x==?20'b1?1??11???1??????11?) z |= 4'b1000; 
	if(x==?20'b?1??011???????0?111?) z |= 4'b1100; 
	if(x==?20'b1???111?????????111?) z |= 4'b1000; 
	if(x==?20'b?????1?1?????1?1?1?1) z |= 4'b1001; 
	if(x==?20'b111?????1????????111) z |= 4'b1000; 
	if(x==?20'b?1????1????10???111?) z |= 4'b0100; 
	if(x==?20'b??1??11?1??1????1??1) z |= 4'b0100; 
	if(x==?20'b?1??1?1??1????0??11?) z |= 4'b1000; 
	if(x==?20'b??????11??11????1?1?) z |= 4'b0001; 
	if(x==?20'b??11??1????1????1?11) z |= 4'b0100; 
	if(x==?20'b???1?111????????111?) z |= 4'b0100; 
	if(x==?20'b?11?11??1???????1??1) z |= 4'b1000; 
	if(x==?20'b?1??11???????00?1??1) z |= 4'b1000; 
	if(x==?20'b?1?????1???1??0?11?1) z |= 4'b0100; 
	if(x==?20'b?1??111?1????????11?) z |= 4'b1000; 
	if(x==?20'b??1???11?????00?1??1) z |= 4'b0100; 
	if(x==?20'b?111???????1?????111) z |= 4'b0100; 
	if(x==?20'b??1??1?1??1??0???11?) z |= 4'b0100; 
	if(x==?20'b111?????1???????11?1) z |= 4'b1000; 
	if(x==?20'b?11?11?????1????1??1) z |= 4'b1000; 
	if(x==?20'b????11??1????0??111?) z |= 4'b1000; 
	if(x==?20'b?11???11???1????1??1) z |= 4'b0100; 
	if(x==?20'b111??1???1???????11?) z |= 4'b1000; 
	if(x==?20'b?1??111?1???????11??) z |= 4'b1000; 
	if(x==?20'b?111???????1????11?1) z |= 4'b0100; 
	if(x==?20'b??1??111???1?????11?) z |= 4'b0100; 
	if(x==?20'b?111??1???1??????11?) z |= 4'b0100; 
	if(x==?20'b1?1?11??????????111?) z |= 4'b1000; 
	if(x==?20'b?1?1??11????????111?) z |= 4'b0100; 
	if(x==?20'b??????11???1??0?111?) z |= 4'b0100; 
	if(x==?20'b111??1???1??????11??) z |= 4'b1000; 
	if(x==?20'b???1??1?0???0????1?1) z |= 4'b0100; 
	if(x==?20'b??1??111???1????11??) z |= 4'b0100; 
	if(x==?20'b1?1??1??1???????111?) z |= 4'b1000; 
	if(x==?20'b?111??1???1?????11??) z |= 4'b0100; 
	if(x==?20'b?11?11??1????????11?) z |= 4'b1000; 
	if(x==?20'b1????1?????0???0?1?1) z |= 4'b1000; 
	if(x==?20'b?1???111??1?????1??1) z |= 4'b0100; 
	if(x==?20'b????11???11?????1?1?) z |= 4'b0010; 
	if(x==?20'b??????11?11?????1?1?) z |= 4'b0001; 
	if(x==?20'b?1?1??1????1????111?) z |= 4'b0100; 
	if(x==?20'b?11???11???1?????11?) z |= 4'b0100; 
	if(x==?20'b?1??0?1??????0??111?) z |= 4'b0100; 
	if(x==?20'b??1??1?0??????0?111?) z |= 4'b1000; 
	if(x==?20'b??1?111??1???????11?) z |= 4'b1000; 
	if(x==?20'b??1?11??1???????1?11) z |= 4'b1000; 
	if(x==?20'b?1???111??1??????11?) z |= 4'b0100; 
	if(x==?20'b??1?11?????1????1?11) z |= 4'b1000; 
	if(x==?20'b?1????11???1????1?11) z |= 4'b0100; 
	if(x==?20'b????111?1???????111?) z |= 4'b1000; 
	if(x==?20'b????1?10???0?????1?1) z |= 4'b1000; 
	if(x==?20'b????01?10????????1?1) z |= 4'b0100; 
	if(x==?20'b111??11?????????1??1) z |= 4'b1000; 
	if(x==?20'b?????1???1??1?1??1??) z |= 4'b0010; 
	if(x==?20'b?111?11?????????1??1) z |= 4'b0100; 
	if(x==?20'b?11??1????0?????1?11) z |= 4'b1000; 
	if(x==?20'b??????1???1??1?1?1??) z |= 4'b0001; 
	if(x==?20'b?11???1??0??????1?11) z |= 4'b0100; 
	if(x==?20'b?????111???1????111?) z |= 4'b0100; 
	if(x==?20'b??1?????1????00?11?1) z |= 4'b1000; 
	if(x==?20'b?11?11???????0??1??1) z |= 4'b1000; 
	if(x==?20'b?11?11????????0?1??1) z |= 4'b1000; 
	if(x==?20'b?11???11?????0??1??1) z |= 4'b0100; 
	if(x==?20'b?11???11??????0?1??1) z |= 4'b0100; 
	if(x==?20'b?11?0?1?????????1?11) z |= 4'b0100; 
	if(x==?20'b?11??1?0????????1?11) z |= 4'b1000; 
	if(x==?20'b?1?????????1?00?11?1) z |= 4'b0100; 
	if(x==?20'b??1?11??1???????111?) z |= 4'b1000; 
	if(x==?20'b?11?11????1?????11??) z |= 4'b1000; 
	if(x==?20'b?11???11??1?????11??) z |= 4'b0100; 
	if(x==?20'b?1???110????????111?) z |= 4'b1000; 
	if(x==?20'b??1?011?????????111?) z |= 4'b0100; 
	if(x==?20'b?11??1??1?1?????11??) z |= 4'b1000; 
	if(x==?20'b?1????11???1????111?) z |= 4'b0100; 
	if(x==?20'b?????1??1??0???0?1?1) z |= 4'b1000; 
	if(x==?20'b?????????1???1?1?111) z |= 4'b1000; 
	if(x==?20'b?11???1??1?1????11??) z |= 4'b0100; 
	if(x==?20'b??????1?0??10????1?1) z |= 4'b0100; 
	if(x==?20'b?1?1??1??????0??111?) z |= 4'b0100; 
	if(x==?20'b1?1??1???????0??111?) z |= 4'b1000; 
	if(x==?20'b?1?1??1???????0?111?) z |= 4'b0100; 
	if(x==?20'b?11?11???????0???11?) z |= 4'b1000; 
	if(x==?20'b1?1??1????????0?111?) z |= 4'b1000; 
	if(x==?20'b?1???1??11??????1?11) z |= 4'b1000; 
	if(x==?20'b?11?11????????0??11?) z |= 4'b1000; 
	if(x==?20'b?11???11?????0???11?) z |= 4'b0100; 
	if(x==?20'b??????????1?1?1??111) z |= 4'b0100; 
	if(x==?20'b?11???11??????0??11?) z |= 4'b0100; 
	if(x==?20'b?11?1???1???????111?) z |= 4'b1000; 
	if(x==?20'b?11??11??????00?1??1) z |= 4'b1100; 
	if(x==?20'b?11??1??1????0???11?) z |= 4'b1000; 
	if(x==?20'b?????11??????1?1?1?1) z |= 4'b1000; 
	if(x==?20'b?????11?????1?1??1?1) z |= 4'b0100; 
	if(x==?20'b??1???1???11????1?11) z |= 4'b0100; 
	if(x==?20'b?????11?11??????1?1?) z |= 4'b0010; 
	if(x==?20'b?11????1???1????111?) z |= 4'b0100; 
	if(x==?20'b?11???1????1??0??11?) z |= 4'b0100; 
	if(x==?20'b1???1?1????0?????1?1) z |= 4'b1000; 
	if(x==?20'b?11?????11??????1?11) z |= 4'b0100; 
	if(x==?20'b???1?1?10????????1?1) z |= 4'b0100; 
	if(x==?20'b?????11???11????1?1?) z |= 4'b0001; 
	if(x==?20'b??1?1??1?1???1??11??) z |= 4'b1100; 
	if(x==?20'b?1??1??1?1???1??11??) z |= 4'b1100; 
	if(x==?20'b???1??1??1??1???11??) z |= 4'b0100; 
	if(x==?20'b?????11?????11??1??1) z |= 4'b0110; 
	if(x==?20'b1????1??1??0?????1?1) z |= 4'b1000; 
	if(x==?20'b???1?1???1??1???11??) z |= 4'b0100; 
	if(x==?20'b??1?1??1??1??1??11??) z |= 4'b1100; 
	if(x==?20'b?1??1??1??1??1??11??) z |= 4'b1100; 
	if(x==?20'b?11???????11????1?11) z |= 4'b1000; 
	if(x==?20'b???1??1?0??1?????1?1) z |= 4'b0100; 
	if(x==?20'b?????????1??1?1??11?) z |= 4'b0010; 
	if(x==?20'b?111??1?????????1?11) z |= 4'b0100; 
	if(x==?20'b???1?1????1?1???11??) z |= 4'b0100; 
	if(x==?20'b111??1??????????1?11) z |= 4'b1000; 
	if(x==?20'b??????????1??1?1?11?) z |= 4'b0001; 
	if(x==?20'b1?????1??1?????111??) z |= 4'b1000; 
	if(x==?20'b??1?1??1?1????1?11??) z |= 4'b1100; 
	if(x==?20'b?1??1??1?1????1?11??) z |= 4'b1100; 
	if(x==?20'b1?????1???1????111??) z |= 4'b1000; 
	if(x==?20'b??1?1??1??1???1?11??) z |= 4'b1100; 
	if(x==?20'b?11?????1????0??11?1) z |= 4'b1000; 
	if(x==?20'b?1??1??1??1???1?11??) z |= 4'b1100; 
	if(x==?20'b1????1????1????111??) z |= 4'b1000; 
	if(x==?20'b1???11?????????0?1?1) z |= 4'b1000; 
	if(x==?20'b?11?111??????????11?) z |= 4'b1000; 
	if(x==?20'b???1??11????0????1?1) z |= 4'b0100; 
	if(x==?20'b?????11???????111??1) z |= 4'b1001; 
	if(x==?20'b?11??111?????????11?) z |= 4'b0100; 
	if(x==?20'b?11????????1??0?11?1) z |= 4'b0100; 
	if(x==?20'b??1?11???????0??111?) z |= 4'b1000; 
	if(x==?20'b?1????11??????0?111?) z |= 4'b0100; 
	if(x==?20'b??????1?0???0?0??1?1) z |= 4'b0100; 
	if(x==?20'b??1??1??1????0??111?) z |= 4'b1000; 
	if(x==?20'b??1??1??1?????0?111?) z |= 4'b1000; 
	if(x==?20'b?????1?????0?0?0?1?1) z |= 4'b1000; 
	if(x==?20'b??????1??????1?1?1?1) z |= 4'b0001; 
	if(x==?20'b?1????1????1?0??111?) z |= 4'b0100; 
	if(x==?20'b?1????1????1??0?111?) z |= 4'b0100; 
	if(x==?20'b?????1??????1?1??1?1) z |= 4'b0010; 
	if(x==?20'b?????1???????1?1?111) z |= 4'b1000; 
	if(x==?20'b??????1?????1?1??111) z |= 4'b0100; 
	if(x==?20'b????1?1?1??0?????1?1) z |= 4'b1000; 
	if(x==?20'b?11?11??????????1?11) z |= 4'b0100; 
	if(x==?20'b?11???11????????1?11) z |= 4'b1000; 
	if(x==?20'b?????1?10??1?????1?1) z |= 4'b0100; 
	if(x==?20'b?1???????????1?1?111) z |= 4'b1000; 
	if(x==?20'b??1?????????1?1??111) z |= 4'b0100; 
	if(x==?20'b???1??1?0?????0??1?1) z |= 4'b0100; 
	if(x==?20'b?11??1??1???????1?11) z |= 4'b1000; 
	if(x==?20'b1????1?????0?0???1?1) z |= 4'b1000; 
	if(x==?20'b??1?111?????????111?) z |= 4'b1000; 
	if(x==?20'b????1???1???1???11??) z |= 4'b0010; 
	if(x==?20'b?11???1????1????1?11) z |= 4'b0100; 
	if(x==?20'b?1???111????????111?) z |= 4'b0100; 
	if(x==?20'b????11??1??????0?1?1) z |= 4'b1000; 
	if(x==?20'b??????11???10????1?1) z |= 4'b0100; 
	if(x==?20'b1?????1??1???1??11??) z |= 4'b1000; 
	if(x==?20'b???1??1??1???1??11??) z |= 4'b0100; 
	if(x==?20'b???1?1???1???1??11??) z |= 4'b0100; 
	if(x==?20'b???????1???1???111??) z |= 4'b0001; 
	if(x==?20'b1?????1???1??1??11??) z |= 4'b1000; 
	if(x==?20'b1????1????1??1??11??) z |= 4'b1000; 
	if(x==?20'b??1??1??1??1?1??11??) z |= 4'b1100; 
	if(x==?20'b???1?1????1??1??11??) z |= 4'b0100; 
	if(x==?20'b?1????1?0???0????1?1) z |= 4'b0100; 
	if(x==?20'b1?????1??1????1?11??) z |= 4'b1000; 
	if(x==?20'b???1??1??1????1?11??) z |= 4'b0100; 
	if(x==?20'b??1??1?????0???0?1?1) z |= 4'b1000; 
	if(x==?20'b???1?1???1????1?11??) z |= 4'b0100; 
	if(x==?20'b?????????????1?1?111) z |= 4'b0001; 
	if(x==?20'b1?????1???1???1?11??) z |= 4'b1000; 
	if(x==?20'b????????????1?1??111) z |= 4'b0010; 
	if(x==?20'b1????1????1???1?11??) z |= 4'b1000; 
	if(x==?20'b??1??1??1??1??1?11??) z |= 4'b1100; 
	if(x==?20'b???1?1????1???1?11??) z |= 4'b0100; 
	if(x==?20'b????????????11??1?11) z |= 4'b0010; 
	if(x==?20'b1???11??1????????1?1) z |= 4'b1000; 
	if(x==?20'b?11?????0??0?????111) z |= 4'b1100; 
	if(x==?20'b????1????1??1???11??) z |= 4'b0010; 
	if(x==?20'b???????1?1??1???111?) z |= 4'b0100; 
	if(x==?20'b1????110?????????1?1) z |= 4'b1000; 
	if(x==?20'b???1011??????????1?1) z |= 4'b0100; 
	if(x==?20'b???1??11???1?????1?1) z |= 4'b0100; 
	if(x==?20'b???????1??1?1???111?) z |= 4'b0100; 
	if(x==?20'b?1??111???0????????1) z |= 4'b1000; 
	if(x==?20'b???????1?1?????111??) z |= 4'b0001; 
	if(x==?20'b????1????1?????1111?) z |= 4'b1000; 
	if(x==?20'b??????????????111?11) z |= 4'b0001; 
	if(x==?20'b????1?1??1???1???1??) z |= 4'b0010; 
	if(x==?20'b?????1??1??0?0???1?1) z |= 4'b1000; 
	if(x==?20'b???????1??1????111??) z |= 4'b0001; 
	if(x==?20'b????1?????1????1111?) z |= 4'b1000; 
	if(x==?20'b??1??111?0?????????1) z |= 4'b0100; 
	if(x==?20'b?1?1??1?0????????1?1) z |= 4'b0100; 
	if(x==?20'b??????1?0??1??0??1?1) z |= 4'b0100; 
	if(x==?20'b1?1??1?????0?????1?1) z |= 4'b1000; 
	if(x==?20'b?????1??1?1??1???1??) z |= 4'b0010; 
	if(x==?20'b??1?0???0????????111) z |= 4'b0100; 
	if(x==?20'b?11??????????11?1?11) z |= 4'b1100; 
	if(x==?20'b??????1?1?1??1???11?) z |= 4'b0100; 
	if(x==?20'b?1?????0???0?????111) z |= 4'b1000; 
	if(x==?20'b??1????011???????111) z |= 4'b1100; 
	if(x==?20'b?????1?1??1???1??1??) z |= 4'b0001; 
	if(x==?20'b??????1??1?1?1???11?) z |= 4'b0100; 
	if(x==?20'b??????1??1?1??1??1??) z |= 4'b0001; 
	if(x==?20'b??1???1?1???1???11??) z |= 4'b0100; 
	if(x==?20'b?????1??1?1???1??11?) z |= 4'b1000; 
	if(x==?20'b?1??0?????11?????111) z |= 4'b1100; 
	if(x==?20'b??11??1?????0????1?1) z |= 4'b0100; 
	if(x==?20'b11???1?????????0?1?1) z |= 4'b1000; 
	if(x==?20'b?????1???1?1??1??11?) z |= 4'b1000; 
	if(x==?20'b????1???1????1??11??) z |= 4'b0010; 
	if(x==?20'b????1??0?1???????111) z |= 4'b1000; 
	if(x==?20'b????0??1??1??????111) z |= 4'b0100; 
	if(x==?20'b???????1???1?1??11??) z |= 4'b0001; 
	if(x==?20'b????1???1?????1?11??) z |= 4'b0010; 
	if(x==?20'b?1???1?????1???111??) z |= 4'b1000; 
	if(x==?20'b1???11???????0???1?1) z |= 4'b1000; 
	if(x==?20'b1???11????????0??1?1) z |= 4'b1000; 
	if(x==?20'b???1??11?????0???1?1) z |= 4'b0100; 
	if(x==?20'b???1??11??????0??1?1) z |= 4'b0100; 
	if(x==?20'b???????1???1??1?11??) z |= 4'b0001; 
	if(x==?20'b1?1?????1?1??????1?1) z |= 4'b1000; 
	if(x==?20'b?1?1????1?1??????1?1) z |= 4'b0100; 
	if(x==?20'b??????1??11??1???11?) z |= 4'b0100; 
	if(x==?20'b1??????11???????11?1) z |= 4'b1000; 
	if(x==?20'b??1?1?1????0?????1?1) z |= 4'b1000; 
	if(x==?20'b1?1??????1?1?????1?1) z |= 4'b1000; 
	if(x==?20'b?1??1?1????0?????1?1) z |= 4'b1000; 
	if(x==?20'b?1?1?????1?1?????1?1) z |= 4'b0100; 
	if(x==?20'b1????1??1?????0??1?1) z |= 4'b1000; 
	if(x==?20'b??1??1?10????????1?1) z |= 4'b0100; 
	if(x==?20'b?1???1?10????????1?1) z |= 4'b0100; 
	if(x==?20'b???11??????1????11?1) z |= 4'b0100; 
	if(x==?20'b1?????10????????11?1) z |= 4'b1000; 
	if(x==?20'b?1??1?10?????????1?1) z |= 4'b1000; 
	if(x==?20'b???1??1????1?0???1?1) z |= 4'b0100; 
	if(x==?20'b???101??????????11?1) z |= 4'b0100; 
	if(x==?20'b??11????0????????111) z |= 4'b0100; 
	if(x==?20'b?1????1??1??1???11??) z |= 4'b0100; 
	if(x==?20'b?????1??1???1???11??) z |= 4'b0010; 
	if(x==?20'b??1??1??1??0?????1?1) z |= 4'b1000; 
	if(x==?20'b?????1???11???1??11?) z |= 4'b1000; 
	if(x==?20'b??1??1???1??1???11??) z |= 4'b0100; 
	if(x==?20'b?1???1???1??1???11??) z |= 4'b0100; 
	if(x==?20'b??1?01?1?????????1?1) z |= 4'b0100; 
	if(x==?20'b11?????????0?????111) z |= 4'b1000; 
	if(x==?20'b1???????1??1????11?1) z |= 4'b1000; 
	if(x==?20'b?1?1?????????1???111) z |= 4'b0100; 
	if(x==?20'b???1????1??1????11?1) z |= 4'b0100; 
	if(x==?20'b?1????1?0??1?????1?1) z |= 4'b0100; 
	if(x==?20'b??1??1????1?1???11??) z |= 4'b0100; 
	if(x==?20'b?1???1????1?1???11??) z |= 4'b0100; 
	if(x==?20'b????1????1???1??11??) z |= 4'b0010; 
	if(x==?20'b??1???1??1?????111??) z |= 4'b1000; 
	if(x==?20'b?1????1??1?????111??) z |= 4'b1000; 
	if(x==?20'b????????1?1??1???11?) z |= 4'b0010; 
	if(x==?20'b????1????1???1??111?) z |= 4'b1000; 
	if(x==?20'b????1?????1??1??11??) z |= 4'b0010; 
	if(x==?20'b??1???1???1????111??) z |= 4'b1000; 
	if(x==?20'b?1????1???1????111??) z |= 4'b1000; 
	if(x==?20'b???????1??1??1??11??) z |= 4'b0001; 
	if(x==?20'b???????1?1???1??111?) z |= 4'b0100; 
	if(x==?20'b????1?????1??1??111?) z |= 4'b1000; 
	if(x==?20'b??1??1????1????111??) z |= 4'b1000; 
	if(x==?20'b1?1???????????1??111) z |= 4'b1000; 
	if(x==?20'b??????1????1???111??) z |= 4'b0001; 
	if(x==?20'b??1?11?????????0?1?1) z |= 4'b1000; 
	if(x==?20'b????1???????1???11?1) z |= 4'b0010; 
	if(x==?20'b???????1??1??1??111?) z |= 4'b0100; 
	if(x==?20'b????1????1????1?11??) z |= 4'b0010; 
	if(x==?20'b?1????11????0????1?1) z |= 4'b0100; 
	if(x==?20'b1???1????1???????111) z |= 4'b1000; 
	if(x==?20'b???????1?1????1?11??) z |= 4'b0001; 
	if(x==?20'b????1????1????1?111?) z |= 4'b1000; 
	if(x==?20'b????1?????1???1?11??) z |= 4'b0010; 
	if(x==?20'b????1?????????0011?1) z |= 4'b1000; 
	if(x==?20'b?????????1?1??1??11?) z |= 4'b0001; 
	if(x==?20'b????1?1??1?1?????1?1) z |= 4'b1000; 
	if(x==?20'b???????1????00??11?1) z |= 4'b0100; 
	if(x==?20'b???????1??1???1?11??) z |= 4'b0001; 
	if(x==?20'b???????1?1????1?111?) z |= 4'b0100; 
	if(x==?20'b?1???1??1??????0?1?1) z |= 4'b1000; 
	if(x==?20'b????1?????1???1?111?) z |= 4'b1000; 
	if(x==?20'b?????1?11?1??????1?1) z |= 4'b0100; 
	if(x==?20'b???1???1??1??????111) z |= 4'b0100; 
	if(x==?20'b?????????????11?1?11) z |= 4'b0011; 
	if(x==?20'b1?1??????11??????1?1) z |= 4'b1000; 
	if(x==?20'b???????1??1???1?111?) z |= 4'b0100; 
	if(x==?20'b?1?1?????11??????1?1) z |= 4'b0100; 
	if(x==?20'b???????1???????111?1) z |= 4'b0001; 
	if(x==?20'b??1???1????10????1?1) z |= 4'b0100; 
	if(x==?20'b??????1111??????1??1) z |= 4'b0100; 
	if(x==?20'b??????1??1??1???11??) z |= 4'b0010; 
	if(x==?20'b?????1???1??1???11??) z |= 4'b0010; 
	if(x==?20'b11???????11?????1??1) z |= 4'b1000; 
	if(x==?20'b??11?????11?????1??1) z |= 4'b0100; 
	if(x==?20'b????11????11????1??1) z |= 4'b1000; 
	if(x==?20'b?????1????1?1???11??) z |= 4'b0010; 
	if(x==?20'b????11??1????0???1?1) z |= 4'b1000; 
	if(x==?20'b????11??1?????0??1?1) z |= 4'b1000; 
	if(x==?20'b?1????10?1???????1?1) z |= 4'b1000; 
	if(x==?20'b??1??1????1??1???1?1) z |= 4'b0100; 
	if(x==?20'b??????1??1?????111??) z |= 4'b0001; 
	if(x==?20'b??1???1?1????1??11??) z |= 4'b0100; 
	if(x==?20'b11??1?1??????????1?1) z |= 4'b1000; 
	if(x==?20'b1?1?11???????????1?1) z |= 4'b1000; 
	if(x==?20'b??1?01????1??????1?1) z |= 4'b0100; 
	if(x==?20'b?1????1??1????1??1?1) z |= 4'b1000; 
	if(x==?20'b??????1???1????111??) z |= 4'b0001; 
	if(x==?20'b?1?1??11?????????1?1) z |= 4'b0100; 
	if(x==?20'b?????1????1????111??) z |= 4'b0001; 
	if(x==?20'b??????11???1?0???1?1) z |= 4'b0100; 
	if(x==?20'b??11?1?1?????????1?1) z |= 4'b0100; 
	if(x==?20'b??????11???1??0??1?1) z |= 4'b0100; 
	if(x==?20'b?1??1??????0?????111) z |= 4'b1000; 
	if(x==?20'b??1????10????????111) z |= 4'b0100; 
	if(x==?20'b1???1?????????0?11?1) z |= 4'b1000; 
	if(x==?20'b???1???1?????0??11?1) z |= 4'b0100; 
	if(x==?20'b11???1??1????????1?1) z |= 4'b1000; 
	if(x==?20'b?1??1??0?????????111) z |= 4'b1000; 
	if(x==?20'b????????1???1???111?) z |= 4'b0010; 
	if(x==?20'b?1??????1??0?????111) z |= 4'b1000; 
	if(x==?20'b??1?0??1?????????111) z |= 4'b0100; 
	if(x==?20'b?1????1?0?????0??1?1) z |= 4'b0100; 
	if(x==?20'b??11??1????1?????1?1) z |= 4'b0100; 
	if(x==?20'b??1??1?????0?0???1?1) z |= 4'b1000; 
	if(x==?20'b?1???1?????1??1?11??) z |= 4'b1000; 
	if(x==?20'b??1?????0??1?????111) z |= 4'b0100; 
	if(x==?20'b????11???11?????1??1) z |= 4'b1000; 
	if(x==?20'b??????11?11?????1??1) z |= 4'b0100; 
	if(x==?20'b??1???1??1???1???11?) z |= 4'b0100; 
	if(x==?20'b???????????1???1111?) z |= 4'b0001; 
	if(x==?20'b????1???11???????111) z |= 4'b1000; 
	if(x==?20'b?1???1???10?????11??) z |= 4'b1000; 
	if(x==?20'b??1???1??1???1??11??) z |= 4'b1000; 
	if(x==?20'b?1??1??????????011?1) z |= 4'b1000; 
	if(x==?20'b??1???1??01?????11??) z |= 4'b0100; 
	if(x==?20'b?????1??1????1??11??) z |= 4'b0010; 
	if(x==?20'b??1??1???1???1??11??) z |= 4'b0100; 
	if(x==?20'b?1???1???1???1??11??) z |= 4'b0100; 
	if(x==?20'b??1????1????0???11?1) z |= 4'b0100; 
	if(x==?20'b??1???1?????0?0??1?1) z |= 4'b0100; 
	if(x==?20'b?1???1???????0?0?1?1) z |= 4'b1000; 
	if(x==?20'b??1???1???1??1??11??) z |= 4'b1000; 
	if(x==?20'b?1????1???1??1??11??) z |= 4'b1000; 
	if(x==?20'b???????1??11?????111) z |= 4'b0100; 
	if(x==?20'b?1???1????1???1??11?) z |= 4'b1000; 
	if(x==?20'b??????1????1?1??11??) z |= 4'b0001; 
	if(x==?20'b11????1??1???????1?1) z |= 4'b1000; 
	if(x==?20'b?????1??1?????1?11??) z |= 4'b0010; 
	if(x==?20'b??1??1???1????1?11??) z |= 4'b0100; 
	if(x==?20'b?1???1???1????1?11??) z |= 4'b0100; 
	if(x==?20'b?????????1??1???111?) z |= 4'b0010; 
	if(x==?20'b??1???1???1???1?11??) z |= 4'b1000; 
	if(x==?20'b??11?1????1??????1?1) z |= 4'b0100; 
	if(x==?20'b?1????1???1???1?11??) z |= 4'b1000; 
	if(x==?20'b?1??1????1????0??1?1) z |= 4'b1000; 
	if(x==?20'b?1???1????1???1?11??) z |= 4'b0100; 
	if(x==?20'b????1????????1??11?1) z |= 4'b0010; 
	if(x==?20'b??????1????1??1?11??) z |= 4'b0001; 
	if(x==?20'b???????1?????1??11?1) z |= 4'b0001; 
	if(x==?20'b?1??1?1?1????????1?1) z |= 4'b1000; 
	if(x==?20'b??1????1??1??0???1?1) z |= 4'b0100; 
	if(x==?20'b??1?11??1????????1?1) z |= 4'b1000; 
	if(x==?20'b11??1????????????111) z |= 4'b1000; 
	if(x==?20'b??????????1????1111?) z |= 4'b0001; 
	if(x==?20'b??11???1?????????111) z |= 4'b0100; 
	if(x==?20'b????1?????????1?11?1) z |= 4'b0010; 
	if(x==?20'b????1???1?????0?11?1) z |= 4'b1000; 
	if(x==?20'b???????1??????1?11?1) z |= 4'b0001; 
	if(x==?20'b??1??110?????????1?1) z |= 4'b1000; 
	if(x==?20'b?1??011??????????1?1) z |= 4'b0100; 
	if(x==?20'b?1????11???1?????1?1) z |= 4'b0100; 
	if(x==?20'b??1??1?1???1?????1?1) z |= 4'b0100; 
	if(x==?20'b11??1???????????11?1) z |= 4'b1000; 
	if(x==?20'b?1?1??1??????0???1?1) z |= 4'b0100; 
	if(x==?20'b11???1???????0???1?1) z |= 4'b1000; 
	if(x==?20'b??11???1????????11?1) z |= 4'b0100; 
	if(x==?20'b??11??1???????0??1?1) z |= 4'b0100; 
	if(x==?20'b1?1??1????????0??1?1) z |= 4'b1000; 
	if(x==?20'b???????1???1?0??11?1) z |= 4'b0100; 
	if(x==?20'b?????1???1???1??11??) z |= 4'b0001; 
	if(x==?20'b??????1?????0?0??111) z |= 4'b0100; 
	if(x==?20'b?????1???????0?0?111) z |= 4'b1000; 
	if(x==?20'b??????1?????1???11?1) z |= 4'b0010; 
	if(x==?20'b??????1??1???1??11??) z |= 4'b0011; 
	if(x==?20'b??????1???1???1?11??) z |= 4'b0010; 
	if(x==?20'b?11?1??1?????????111) z |= 4'b1100; 
	if(x==?20'b??????1???1??1??11??) z |= 4'b0011; 
	if(x==?20'b?????1????1??1??11??) z |= 4'b0011; 
	if(x==?20'b???1??1?1???????111?) z |= 4'b0100; 
	if(x==?20'b?????1?????????111?1) z |= 4'b0001; 
	if(x==?20'b???1?1??1???????111?) z |= 4'b0100; 
	if(x==?20'b????????1????1??111?) z |= 4'b0010; 
	if(x==?20'b??????1??1????1?11??) z |= 4'b0011; 
	if(x==?20'b?????11?11??????1??1) z |= 4'b0100; 
	if(x==?20'b?????1???1????1?11??) z |= 4'b0011; 
	if(x==?20'b1?????1????1????111?) z |= 4'b1000; 
	if(x==?20'b1????1?????1????111?) z |= 4'b1000; 
	if(x==?20'b?11???1?????0????1?1) z |= 4'b0100; 
	if(x==?20'b?1????1?11???????1?1) z |= 4'b1000; 
	if(x==?20'b?????1????1???1?11??) z |= 4'b0011; 
	if(x==?20'b?11??1?????????0?1?1) z |= 4'b1000; 
	if(x==?20'b???????????1?1??111?) z |= 4'b0001; 
	if(x==?20'b?1?1?????1???????111) z |= 4'b0100; 
	if(x==?20'b????????1?????1?111?) z |= 4'b0010; 
	if(x==?20'b1?1???????1??????111) z |= 4'b1000; 
	if(x==?20'b?????11???11????1??1) z |= 4'b1000; 
	if(x==?20'b???????????1??1?111?) z |= 4'b0001; 
	if(x==?20'b??1??1????11?????1?1) z |= 4'b0100; 
	if(x==?20'b?1??1???1????????111) z |= 4'b1000; 
	if(x==?20'b??1?11???????0???1?1) z |= 4'b1000; 
	if(x==?20'b??1?11????????0??1?1) z |= 4'b1000; 
	if(x==?20'b?1????11?????0???1?1) z |= 4'b0100; 
	if(x==?20'b?1????11??????0??1?1) z |= 4'b0100; 
	if(x==?20'b?1??1???1???????11?1) z |= 4'b1000; 
	if(x==?20'b????1????????00?11?1) z |= 4'b1000; 
	if(x==?20'b??1????1???1?????111) z |= 4'b0100; 
	if(x==?20'b??1????11???????11?1) z |= 4'b1000; 
	if(x==?20'b?1?????11???????11?1) z |= 4'b1000; 
	if(x==?20'b?1???1??1????0???1?1) z |= 4'b1000; 
	if(x==?20'b???????1?????00?11?1) z |= 4'b0100; 
	if(x==?20'b??1??1??1?????0??1?1) z |= 4'b1000; 
	if(x==?20'b?1??11???1???????11?) z |= 4'b1000; 
	if(x==?20'b?????????1???1??111?) z |= 4'b0001; 
	if(x==?20'b??1?1??????1????11?1) z |= 4'b0100; 
	if(x==?20'b??1???11?1???????11?) z |= 4'b0100; 
	if(x==?20'b?1??1??????1????11?1) z |= 4'b0100; 
	if(x==?20'b??1???10????????11?1) z |= 4'b1000; 
	if(x==?20'b?111??1??????????1?1) z |= 4'b0100; 
	if(x==?20'b?1??1?1???1??????11?) z |= 4'b1000; 
	if(x==?20'b??1??1?1?1???????11?) z |= 4'b0100; 
	if(x==?20'b111??1???????????1?1) z |= 4'b1000; 
	if(x==?20'b?1????1????1?0???1?1) z |= 4'b0100; 
	if(x==?20'b?1??11????1??????11?) z |= 4'b1000; 
	if(x==?20'b?1??01??????????11?1) z |= 4'b0100; 
	if(x==?20'b??1????1???1????11?1) z |= 4'b0100; 
	if(x==?20'b??1???1????1??0??1?1) z |= 4'b0100; 
	if(x==?20'b??1???11??1??????11?) z |= 4'b0100; 
	if(x==?20'b????????????1???1111) z |= 4'b0010; 
	if(x==?20'b??????????1???1?111?) z |= 4'b0010; 
	if(x==?20'b??????????1??1??111?) z |= 4'b0011; 
	if(x==?20'b???????????????11111) z |= 4'b0001; 
	if(x==?20'b?????????1????1?111?) z |= 4'b0011; 
	if(x==?20'b?11??11?1???????1??1) z |= 4'b1100; 
	if(x==?20'b????1?1??1???????11?) z |= 4'b0010; 
	if(x==?20'b?11??11????1????1??1) z |= 4'b1100; 
	if(x==?20'b1?1???1??????????111) z |= 4'b1000; 
	if(x==?20'b?????1?1??1??????11?) z |= 4'b0001; 
	if(x==?20'b?1?1?1???????????111) z |= 4'b0100; 
	if(x==?20'b?????1??1?1??????11?) z |= 4'b0010; 
	if(x==?20'b??????1??1?1?????11?) z |= 4'b0001; 
	if(x==?20'b1?1???1?????????11?1) z |= 4'b1000; 
	if(x==?20'b?11?1?1??????????1?1) z |= 4'b1000; 
	if(x==?20'b?1?1?1??????????11?1) z |= 4'b0100; 
	if(x==?20'b??1???1?????0???111?) z |= 4'b0100; 
	if(x==?20'b?11??1?1?????????1?1) z |= 4'b0100; 
	if(x==?20'b?1???1?????????0111?) z |= 4'b1000; 
	if(x==?20'b?1??1????????0??11?1) z |= 4'b1000; 
	if(x==?20'b??1?1?????????0?11?1) z |= 4'b1000; 
	if(x==?20'b?1??1?????????0?11?1) z |= 4'b1000; 
	if(x==?20'b??1????1?????0??11?1) z |= 4'b0100; 
	if(x==?20'b?1?????1?????0??11?1) z |= 4'b0100; 
	if(x==?20'b?11??1??1????????1?1) z |= 4'b1000; 
	if(x==?20'b??1????1??????0?11?1) z |= 4'b0100; 
	if(x==?20'b?1??????1?????0?11?1) z |= 4'b1000; 
	if(x==?20'b?11???1????1?????1?1) z |= 4'b0100; 
	if(x==?20'b??1????????1?0??11?1) z |= 4'b0100; 
	if(x==?20'b????111???????????11) z |= 4'b0010; 
	if(x==?20'b???????1???1????111?) z |= 4'b0001; 
	if(x==?20'b?????111??????????11) z |= 4'b0001; 
	if(x==?20'b??11??1?????????111?) z |= 4'b0100; 
	if(x==?20'b11???1??????????111?) z |= 4'b1000; 
	if(x==?20'b?????????????1??1111) z |= 4'b0001; 
	if(x==?20'b?11???1??1???????1?1) z |= 4'b1000; 
	if(x==?20'b?11??1????1??????1?1) z |= 4'b0100; 
	if(x==?20'b????1????1??????111?) z |= 4'b0010; 
	if(x==?20'b??????????????1?1111) z |= 4'b0010; 
	if(x==?20'b?1??11??????????1?11) z |= 4'b1000; 
	if(x==?20'b????1?????1?????111?) z |= 4'b0010; 
	if(x==?20'b??1???11????????1?11) z |= 4'b0100; 
	if(x==?20'b???????1??1?????111?) z |= 4'b0001; 
	if(x==?20'b?11?1???????????11?1) z |= 4'b1000; 
	if(x==?20'b?11??1???????0???1?1) z |= 4'b1000; 
	if(x==?20'b?11????1????????11?1) z |= 4'b0100; 
	if(x==?20'b?11???1???????0??1?1) z |= 4'b0100; 
	if(x==?20'b?????11??????11?1??1) z |= 4'b1111; 
	if(x==?20'b?1??11??????????111?) z |= 4'b1000; 
	if(x==?20'b??1???11????????111?) z |= 4'b0100; 
	if(x==?20'b????11??????????1?11) z |= 4'b0010; 
	if(x==?20'b?1????1?1???????111?) z |= 4'b0100; 
	if(x==?20'b??????11????????1?11) z |= 4'b0001; 
	if(x==?20'b??1??1??1???????111?) z |= 4'b0100; 
	if(x==?20'b?1????1????1????111?) z |= 4'b1000; 
	if(x==?20'b??1??1?????1????111?) z |= 4'b1000; 
	if(x==?20'b????????1111??????11) z |= 4'b1100; 
	if(x==?20'b?1???1???????0??111?) z |= 4'b1000; 
	if(x==?20'b??1???1???????0?111?) z |= 4'b0100; 
	if(x==?20'b??????110????????1?1) z |= 4'b0100; 
	if(x==?20'b????11?????0?????1?1) z |= 4'b1000; 
	if(x==?20'b?????1?1?????1???1?1) z |= 4'b0100; 
	if(x==?20'b????1?1???????1??1?1) z |= 4'b1000; 
	if(x==?20'b????1?1??????1???1?1) z |= 4'b0110; 
	if(x==?20'b?????1?1??????1??1?1) z |= 4'b1001; 
	if(x==?20'b??????101???????11?1) z |= 4'b1100; 
	if(x==?20'b????1?1??1?1?????11?) z |= 4'b1100; 
	if(x==?20'b?11???1?????????111?) z |= 4'b0100; 
	if(x==?20'b?????1?11?1??????11?) z |= 4'b1100; 
	if(x==?20'b?11??1??????????111?) z |= 4'b1000; 
	if(x==?20'b????01?????1????11?1) z |= 4'b1100; 
	if(x==?20'b????1?1?1?1??????11?) z |= 4'b1110; 
	if(x==?20'b?????1?1?1?1?????11?) z |= 4'b1101; 
	if(x==?20'b??????1?0????0???1?1) z |= 4'b0100; 
	if(x==?20'b?1????1??1???1??11??) z |= 4'b1100; 
	if(x==?20'b????1111??????????11) z |= 4'b1100; 
	if(x==?20'b?????1?????0??0??1?1) z |= 4'b1000; 
	if(x==?20'b??1??1????1??1??11??) z |= 4'b1100; 
	if(x==?20'b?1???1????1??1??11??) z |= 4'b1100; 
	if(x==?20'b????1?1??11??????11?) z |= 4'b1100; 
	if(x==?20'b??1???1??1????1?11??) z |= 4'b1100; 
	if(x==?20'b?1????1??1????1?11??) z |= 4'b1100; 
	if(x==?20'b?????1???1???1???1??) z |= 4'b0010; 
	if(x==?20'b?????1?1?11??????11?) z |= 4'b1100; 
	if(x==?20'b??1??1????1???1?11??) z |= 4'b1100; 
	if(x==?20'b??????1?????????1111) z |= 4'b0010; 
	if(x==?20'b?????1??????????1111) z |= 4'b0001; 
	if(x==?20'b??????1???1???1??1??) z |= 4'b0001; 
	if(x==?20'b????????111????????1) z |= 4'b0010; 
	if(x==?20'b????1??1?1??????111?) z |= 4'b1100; 
	if(x==?20'b?????????111???????1) z |= 4'b0001; 
	if(x==?20'b????1??1??1?????111?) z |= 4'b1100; 
	if(x==?20'b??????????1??1???111) z |= 4'b0100; 
	if(x==?20'b?????1??????1???11?1) z |= 4'b0110; 
	if(x==?20'b?????????1????1??111) z |= 4'b1000; 
	if(x==?20'b?????11??????1???1?1) z |= 4'b0100; 
	if(x==?20'b??????1????????111?1) z |= 4'b1001; 
	if(x==?20'b?????11???????1??1?1) z |= 4'b1000; 
	if(x==?20'b??1???1?0????????1?1) z |= 4'b0100; 
	if(x==?20'b?1???1?????0?????1?1) z |= 4'b1000; 
	if(x==?20'b?????????1???1???11?) z |= 4'b0010; 
	if(x==?20'b??????????1???1??11?) z |= 4'b0001; 
	if(x==?20'b????1?1???1??????1?1) z |= 4'b1000; 
	if(x==?20'b?????1?1?1???????1?1) z |= 4'b0100; 
	if(x==?20'b?????11?1?1??????11?) z |= 4'b1100; 
	if(x==?20'b?????11??1?1?????11?) z |= 4'b1100; 
	if(x==?20'b??????1?1?1??????1?1) z |= 4'b0100; 
	if(x==?20'b?????1???1?1?????1?1) z |= 4'b1000; 
	if(x==?20'b1????????1??????11?1) z |= 4'b1000; 
	if(x==?20'b???1?????1??????11?1) z |= 4'b0100; 
	if(x==?20'b?????11??11?????1??1) z |= 4'b1100; 
	if(x==?20'b1?????????1?????11?1) z |= 4'b1000; 
	if(x==?20'b??1?????1??1????11?1) z |= 4'b1100; 
	if(x==?20'b?1??????1??1????11?1) z |= 4'b1100; 
	if(x==?20'b???1??????1?????11?1) z |= 4'b0100; 
	if(x==?20'b?????1???????1???1?1) z |= 4'b0010; 
	if(x==?20'b??????1??????1???111) z |= 4'b0100; 
	if(x==?20'b?1??????1?1??????1?1) z |= 4'b1000; 
	if(x==?20'b??1?????1?1??????1?1) z |= 4'b0100; 
	if(x==?20'b??????1???????1??1?1) z |= 4'b0001; 
	if(x==?20'b?1???????1?1?????1?1) z |= 4'b1000; 
	if(x==?20'b???????11???????11?1) z |= 4'b0100; 
	if(x==?20'b??1??????1?1?????1?1) z |= 4'b0100; 
	if(x==?20'b??1?1????1???????111) z |= 4'b1100; 
	if(x==?20'b?????1????????1??111) z |= 4'b1000; 
	if(x==?20'b????1??????1????11?1) z |= 4'b1000; 
	if(x==?20'b??????1?1??1????111?) z |= 4'b1100; 
	if(x==?20'b?????1??1??1????111?) z |= 4'b1100; 
	if(x==?20'b?1?????1??1??????111) z |= 4'b1100; 
	if(x==?20'b?????11??11??????11?) z |= 4'b1100; 
	if(x==?20'b??1??????????1???111) z |= 4'b0100; 
	if(x==?20'b?????1???????1??11?1) z |= 4'b0101; 
	if(x==?20'b?1????????????1??111) z |= 4'b1000; 
	if(x==?20'b??????1???????1?11?1) z |= 4'b1010; 
	if(x==?20'b?11??????11?????1??1) z |= 4'b1100; 
	if(x==?20'b????????1?1??????1?1) z |= 4'b0010; 
	if(x==?20'b?1???????11??????1?1) z |= 4'b1000; 
	if(x==?20'b????1????1??????11?1) z |= 4'b1000; 
	if(x==?20'b??1??????11??????1?1) z |= 4'b0100; 
	if(x==?20'b????111??????????1?1) z |= 4'b1000; 
	if(x==?20'b?????????1?1?????1?1) z |= 4'b0001; 
	if(x==?20'b???????1?1??????11?1) z |= 4'b0100; 
	if(x==?20'b????1?????1?????11?1) z |= 4'b1000; 
	if(x==?20'b?????111?????????1?1) z |= 4'b0100; 
	if(x==?20'b???????1??1?????11?1) z |= 4'b0100; 
	if(x==?20'b????????11??????1??1) z |= 4'b0010; 
	if(x==?20'b???1??1??????????111) z |= 4'b0100; 
	if(x==?20'b1????1???????????111) z |= 4'b1000; 
	if(x==?20'b?????????????1???111) z |= 4'b0010; 
	if(x==?20'b?????11??11?????1?1?) z |= 4'b1111; 
	if(x==?20'b??????????11????1??1) z |= 4'b0001; 
	if(x==?20'b?1??11???????????1?1) z |= 4'b1000; 
	if(x==?20'b??1???11?????????1?1) z |= 4'b0100; 
	if(x==?20'b??????????????1??111) z |= 4'b0001; 
	if(x==?20'b????11???????????111) z |= 4'b1000; 
	if(x==?20'b??????11?????????111) z |= 4'b0100; 
	if(x==?20'b?????????11?????1??1) z |= 4'b0011; 
	if(x==?20'b?????1??1????????111) z |= 4'b1000; 
	if(x==?20'b??????1????1?????111) z |= 4'b0100; 
	if(x==?20'b?????1??1???????11?1) z |= 4'b0100; 
	if(x==?20'b1???????????????1111) z |= 4'b1000; 
	if(x==?20'b???1????????????1111) z |= 4'b0100; 
	if(x==?20'b??????1????1????11?1) z |= 4'b1000; 
	if(x==?20'b??1???1??????0???1?1) z |= 4'b0100; 
	if(x==?20'b?1???1??1???????111?) z |= 4'b1100; 
	if(x==?20'b?1???1????????0??1?1) z |= 4'b1000; 
	if(x==?20'b??1???1????1????111?) z |= 4'b1100; 
	if(x==?20'b??????1??1???????111) z |= 4'b1000; 
	if(x==?20'b?????1????1??????111) z |= 4'b0100; 
	if(x==?20'b??????1??1??????11?1) z |= 4'b1000; 
	if(x==?20'b?????1???1??????11?1) z |= 4'b0100; 
	if(x==?20'b??????1???1?????11?1) z |= 4'b1000; 
	if(x==?20'b?????1????1?????11?1) z |= 4'b0100; 
	if(x==?20'b????????1???????11?1) z |= 4'b0010; 
	if(x==?20'b????????1???????1111) z |= 4'b1000; 
	if(x==?20'b?????1???1???????11?) z |= 4'b0010; 
	if(x==?20'b???????????1????11?1) z |= 4'b0001; 
	if(x==?20'b??????1???1??????11?) z |= 4'b0001; 
	if(x==?20'b????1???????????1111) z |= 4'b1010; 
	if(x==?20'b???????????1????1111) z |= 4'b0100; 
	if(x==?20'b???????1????????1111) z |= 4'b0101; 
	if(x==?20'b?????1???1??????111?) z |= 4'b0101; 
	if(x==?20'b??????1???1?????111?) z |= 4'b1010; 
	if(x==?20'b?????????1??????11?1) z |= 4'b0001; 
	if(x==?20'b??????????1?????11?1) z |= 4'b0010; 
	if(x==?20'b?1????1?????????11?1) z |= 4'b1000; 
	if(x==?20'b??1??1??????????11?1) z |= 4'b0100; 
	if(x==?20'b??????1??????????111) z |= 4'b0001; 
	if(x==?20'b?????1???????????111) z |= 4'b0010; 
	if(x==?20'b????1??1????????11?1) z |= 4'b1100; 
	if(x==?20'b??????1??????1??11?1) z |= 4'b1111; 
	if(x==?20'b???10001111?111?0010) z |= 4'b0100; 
	if(x==?20'b????????1?1??????111) z |= 4'b1100; 
	if(x==?20'b?????1????????1?11?1) z |= 4'b1111; 
	if(x==?20'b?????????1?1?????111) z |= 4'b1100; 
	if(x==?20'b1???1000?111?1110010) z |= 4'b1000; 
	if(x==?20'b?????????11??????111) z |= 4'b1100; 
	if(x==?20'b?????????11?????1?11) z |= 4'b1100; 
	if(x==?20'b????1?1??????????111) z |= 4'b1110; 
	if(x==?20'b?????1?1?????????111) z |= 4'b1101; 
	if(x==?20'b??????1??1???????1?1) z |= 4'b0100; 
	if(x==?20'b?????1????1??????1?1) z |= 4'b1000; 
	if(x==?20'b??1??????1??????11?1) z |= 4'b1100; 
	if(x==?20'b?1???????1??????11?1) z |= 4'b1100; 
	if(x==?20'b??1???????1?????11?1) z |= 4'b1100; 
	if(x==?20'b?1????????1?????11?1) z |= 4'b1100; 
	if(x==?20'b?????????1???????1?1) z |= 4'b0010; 
	if(x==?20'b??????????1??????1?1) z |= 4'b0001; 
	if(x==?20'b?????????1??????1111) z |= 4'b1100; 
	if(x==?20'b?????11??????????111) z |= 4'b1100; 
	if(x==?20'b??????1??1??????111?) z |= 4'b1111; 
	if(x==?20'b??????????1?????1111) z |= 4'b1100; 
	if(x==?20'b?????1????1?????111?) z |= 4'b1111; 
	if(x==?20'b?1??0001111?111?0010) z |= 4'b0100; 
	if(x==?20'b?1????1??????????111) z |= 4'b1100; 
	if(x==?20'b??1??1???????????111) z |= 4'b1100; 
	if(x==?20'b??1?1000?111?1110010) z |= 4'b1000; 
	if(x==?20'b?????11?????????1?11) z |= 4'b1111; 
	if(x==?20'b??1?????????????1111) z |= 4'b1100; 
	if(x==?20'b?1??????????????1111) z |= 4'b1100; 
end 
endmodule