`timescale 1ns/100ps
module seq_reco_tb;
logic [255:0] x1 =   256'b1001010000100100000111110101110101001001010111111111001001111111110111111100101111111001111111111111101111000101111100000001111111111111000010101010001111110111111100111011110000001000011101000100011110101111011111111101011110111001110001111010011111111111;
logic [255:0] y1 =   256'b1111111111111111111111111111111111101111111111111111111111111110111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111111111011111111111111111111111111111111111110001111011111111111111111;
logic [255:0] x1_r = 256'b1001010000100100000111110101110101001001010111111111001001111111110111110110101111111001111111111111101111000101111100000001111111111111000010101010001111110111111100111011110000001000011101000100011110101111011111111101011110111001011001111010011111111111;
logic [255:0] y1_r = 256'b1011111111111111111111111111111111101111111111111111111111111111110111110110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111111111101111111111111111111111111111111111111001011111011111111111111;

logic [255:0] x2 = 256'b1111111111011111111111011110011111110111111111110011110001101100001111111111111111011011111111111111011011111111111111111101111111111011111111111111011111001111111100000011111111111111000111111110011111111111111101111111110000011000111111001100111111111111;
logic [255:0] y2 = 256'b1101000110000001111000000000101111010110000000001010000111100011010100010001010000000000001000000000001010101101011101101000011100010000100000110000001110111010000010000000000000011100001100001000000010111110110000000101101100011111000001101110000110111111;
logic [255:0] x2_r = 256'b1101111111011111111111011110101111110111111111111010110101101010001101111111111111011011111111111111011011111111111111111101111111111011111111111111011111101110111110000001111111111111001101111110011111111111111101111111111000011000101111101100101111111111;
logic [255:0] y2_r = 256'b1101000110000001111000000000101111010110000000001010000101101010011100010001010000000000001000000000001010101101011101101000011100010000100000110000001110101110000010000000000000011100001100001000000010111110110000000101101000011111100001101100100110111111;

logic [255:0] x3 = 256'b1001101101100111111100101101111001110111111111001110000101111100000001101111110110000010101010001111110111010100110011010000001000011001000100011010101101011101101001011100110001100001110010011111111110001010000100100000111110101100101001001010111111110001;
logic [255:0] y3 = 256'b1111111111111111100111111111000001111111111111100011111111101111111111111111111111111100001110011111110111011111111111111111111111111111111101111001111111111111111111101111100111111000111111111111111111111111111111111101111111111111111111111111111111101111;
logic [255:0] x3_r = 256'b1001101101100111110110101101101001111111111111001011000101111100000001101111110110000010001110001111110111010100110011010000001000011001000100011010101101011101101001011100110001100001110010011111111110001010000100100000111110101100101001001010111111110001;
logic [255:0] y3_r = 256'b1011111111111111110110111111100001111111111111001011011111111101111111111111111111111110001110001111110111011111111111111111111111111111111101111010111111111111111111111101110011111001110111111111111111111111111111111101111111111111111111111111111111110111;

logic [255:0] x4 = 256'b0000001111000000000101111010110000000101010000111100111010100110011010000000000001001000000001010101101011101101001011100110001100000110010011110111010000010000000100000011100101100101001001010111110110001001101101100111111000101101110001110111111101001110;
logic [255:0] y4 = 256'b1111111101111111111111111111100111111110000001111111111111100011111111101111111111111111111111111100001100011111100110011111111111111111111111111111111101111001111111111111111111101111100110110000111111111111111111101111111111111101101111111111111111110111;
logic [255:0] x4_r = 256'b0000001111000000000101111010110000000101000001111100111010100110011010000000000001001000000001010101001101111101001011010110001100000110010011110111010000010000000100000011100101100101001001010101111110001001101101100111111000101101110001110111111101001110;
logic [255:0] y4_r = 256'b0111111111011111111111111111110011111111000001111101111111100110111111101111111111111111111111111101001100011101101011010111111111111111111111111111111101111001111111111111111111101111101011010100111110111111111111101111111111111101110111111111111111111110;

logic x, y, clk, rst_n, x_reco_r, y_reco_r;
seq_reco DUT(
    .x(x),
    .y(y),
    .clk(clk),
    .rst_n(rst_n),
    .x_reco_r(x_reco_r),
    .y_reco_r(y_reco_r)
);

function fail(
    string signal,
    bit actual_result,
    bit correct_result
);
    $display("TESTCASE FAILED @ time %4.0f: %s caused failure. Was: %b, Should be: %b", $time, signal, actual_result, correct_result);
    $finish;
endfunction

task reset();
    rst_n = 1; #1;
    rst_n = 0; #1;
    rst_n = 1; #1;
endtask

task test_bs(
    input logic [255:0] x_test, y_test, x_r_test, y_r_test
);
    reset();
    for(int i = 255; i >=0; i--) begin
        //$display("%d", i);
        x = x_test[i];
        y = y_test[i];
        //$display("%d%d", x, y);
        @(posedge clk);
        @(negedge clk);
        //$display("%d%d", x_reco_r, y_reco_r);
        if(x_reco_r != x_r_test[i])
            fail("x", x_reco_r, x_r_test[i]);
        if(y_reco_r != y_r_test[i])
            fail("y", y_reco_r, y_r_test[i]);
    end
    $display("PASSED!");
endtask

always #5 clk = ~clk;

initial begin
    clk = 0; 
    test_bs(x1, y1, x1_r, y1_r);
    test_bs(x2, y2, x2_r, y2_r);
    test_bs(x3, y3, x3_r, y3_r);
    test_bs(x4, y4, x4_r, y4_r);
    $finish;
end
endmodule