`timescale 1ns/10ps
module gb4ed_tb;
    
endmodule