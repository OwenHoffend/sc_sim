
`ifndef RECO_TEST_CASES
`define RECO_TEST_CASES
localparam NUM_DEPTHS = 10;
localparam N = 256;
localparam [255:0] tcs [39:0] = {
256'b0000000000111111111111111101111111111111111111111111110111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111010000111111111111110011111111111111111111111111111111111110001110011111111111111111111111111, 256'b0000000000000000000000000000000000000000000000000000000011000000000000000000000001100000000000000000000011110000000000000000100000000000000100000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 256'b1111111111111111111111111101111111111111111111111111110111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111000001111111111111110011111111111111111111111111111111111110001110011111111111111111111111111, 256'b0000000000000000000000000000000000000000000000000000000011000000000000000000000001100000000000000000000011110000000000000000100000000000000100000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 256'b0000000000000101111110011111101111111101110111110000010000111011001000111111111111111111111011111101110011100011110110111111111110010110001001000001111101111101111011011111111111110010011111111101111111001011111110011111111111111011110001011111000000011111, 256'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001100000000000000000000011110000000000000, 256'b1111111110000101111110011111101111111101110111110000010000111011001000111111111111111111111011111101110011100011110110111111111110010110001001000001111101111101111011011111111111110010011111111101111111001011111110011111111111111011110001011111000000011111, 256'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001100000000000000000000011110000000000000, 256'b0000100010010010110001001100001111101111101111011011111111111110010011111111101111111001011111110011111111111111011110001011111000000011111111111110000101111110011111101111111101110111110000010000111011001000111111111111111111111011111101110011100011110110, 256'b0000100010000000000000000000000001000000000000000000000011100000000000000000000011110000000000100000000011111000000100000000110000000000000110000000000000000000000011000010000000000000000000000000000000000000000000000000001000000000001000000000000000000000, 256'b0111111111110010110001001100001111101111101111011011111111111110010011111111101111111001011111110011111111111111011110001011111000000011111111111110000101111110011111101111111101110111110000010000111011001000111111111111111111111011111101110011100011110110, 256'b0000100010000000000000000000000001000000000000000000000011100000000000000000000011110000000000100000000011111000000100000000110000000000000110000000000000000000000011000010000000000000000000000000000000000000000000000000001000000000001000000000000000000000, 256'b0000001000000000000000000000000100010000000000000000000000001000000000000000000000011100000000000000000000001110000000000100000000011111000000000000000110000000000000110000000000000000000000011000010000000000000000000000000000000000000000000000000001000000, 256'b0000001000001010010111001100011100010100100111111111100010101000001000001111101011011100000010101111111100011110001011001111111001011111000011101111111110011100001011111000000011011111101100011000010100011111101110101001100110100000010000110010001001010101, 256'b0000001000000000000000000000000100010000000000000000000000001000000000000000000000011100000000000000000000001110000000000100000000011111000000000000000110000000000000110000000000000000000000011000010000000000000000000000000000000000000000000000000001000000, 256'b1011010111011010010111001100011000011100100111111111100010100001001000001111101011001010010010101111111100010011011011001111111001011011100011101111111110011100001011111000000011011111101100000101010100011111101110101001100110100000010000110010001000110101, 256'b1101000101000010010000011110010110010100100101011111011000100110110110011111100010110111000111011111111100111000010111100000000110111101011000001010101000111110011101010011001101000000100001100100010001101010110101110110100101110011000110000111001001111011, 256'b1101000101011111111111111110111111111111111111111111111011111110110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111101010011011111111111100111111111111111111111111111111111111101110011001111111111011111111111, 256'b1101000101000010010000011110010110010100100101011111011000100110110110011111100010110111000111011111111100111000010111100000000110111101011000001010101000111110011101010011001101000000100001100100010001101010110101110110100101110011000110000111001001111011, 256'b1111111111111111111111111110111111111111111111111111111011111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111100000111111111111111001111111111111111111111111111111111111000111001111111111101111111111111, 256'b0000000111000010000000000000000111100011000000010001000000000000000000000000001000000100001100100000001100010000100000110000001110011000000000000000000000001100000100000000000000011110010000000100100100011111000000100110000110011111100000110000000111000000, 256'b0000000111000010000000000110101111100011000000010001001110101001100110100000001000000100001100100000011100111011100010111001101110011000000000111101110100011100000100000000011001011110010000010101111101111111000000101110011110011111100000110101111111010011, 256'b0000000111000010000000000000000111100011000000010001000000000000000000000000001000000100001100100000001100010000100000110000001110011000000000000000000000001100000100000000000000011110010000000100100100011111000000100110000110011111100000110000000111000000, 256'b1100000011110000000001011110101100000001010100001111001110101001100110100000000000010010000000010101011010111011010010111001100011000001100100111101110100010100000001000000111001011001010010010101111101100010011011011001111110001011011100011101111111010011, 256'b1010110010100100101011111111000001101111110110000110101010111111110111110111110011110000111110011001000101111011101101011101000111111011111001010001111000000100001100100010001101010110101111101100101001001010111110111101001101101110111101000010010000011111, 256'b1010110011100111101011111111000001101111110110000010101010001111110111110100110011010000001000011001000100011010101101011101000111111011111001010001111000000101111110100010001101010110101111101100101001001010111110111101001101101110111101000010010111011111, 256'b1010110010100100101011111111100100110110111011111110010110111100111111111111100111100010111110000000110111111011000001010101000111111011111010011001101000000100001100100010001101010110101111111100101111011000110000111101001111111111000101000010010000011111, 256'b1111111111001111000101111100000001101111110110000010101010001111110111110100110011010000001000011001000100011010101101011111111001011110110001100001111010011111111110001010000100100000111110101100101001001010111111111001001101101110111111100101101111001111, 256'b0000001111000000000101110011110000000101010000111100111010100010001010000000000001000000000001010101101011101101000011100110000100000110010001110111010000010000000000000011100101100001000000010111110110000000101101100011111000001101110000110111111101000110, 256'b0001111111000000010101110011110000011101010000111100111111100110011111111011111111000111111101011111111111111101100011101110000100011111111111110111010000110011111011111111101101111101000000010111110110000001111111111111111110101111110100111111111101000110, 256'b0000001111000000000101111010110000000101010000111100111010100010001010000000000001000000000001010101101011101101000011100110000100000110010001110111010000010000000000000011100101100001000000010111110110000000101101100011111000001101110000110111111101000110, 256'b1111111100101000010010000011111010111010100100101011111111100100111111111011111110010111111100111111111111110111100010111110000000111111111111100001010111100111111011111111011101111100000100001110100010001111111111111111111110101111011100111000111101001111, 256'b1110111111111011111111110011111111111111111111111111101001111111100111111111111111011111111101111111111111111111011111111111111111111111111111111100111110111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111010001111, 256'b1110111111111011111111110011111111000000111111111111101001111111100111111111111111011111111100000110001111110011001111111111111111111110111111111100111110111111101111111111100111100011011000011111111111111110110111111111111110110111111111111111111010011111, 256'b1111111111110011111111111111111111111111111111111110001110011111110111011111111111111111111111111111111111111101111111111111111111111111110111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111000001111, 256'b1110111111111111110111110011111111000000111111111111110001111111100111111111111111011111111100000110001111110011001111111111111111111110111111111110111100111111101111111111100111100011011000011111111111111110110111111111111110110111111111111111111011111111, 256'b0000011000100001000000100000011100010100000000000000000000011000001000000000000000111010001000001001001000111110000001001100001010101111100001100000001100010000000001100001100000000000000000110100110000000100010000000000000000000000000000000001000011001000, 256'b0100011001110001000001101110111100000100010100011111101110111000101010100000010000111010001000011001011010111110010011011100101010100011100001101101111100010000001001100001101001011001010010110100111111100100011011011001111111001011011100011101111111111001, 256'b0000011000100001000000100000011100110000000000000000000000011000001000000000000000111100100000001001001000111110000001001100001100111111000001100000001110000000000001110000100000000000000000111000110000000100010000000000000000000000000000000001000011001000, 256'b1100001011110000000011011110101100000101010100011111101110101001100110100000010000110010001000110101011010111011010010111001100011000011100100111101110100010100001001000001111001011001010010010101111111100010011011011001111111001011011100011101111111110011
};
`endif
