
`ifndef RECO_TEST_CASES
`define RECO_TEST_CASES
localparam NUM_DEPTHS = 2;
localparam N = 256;
localparam [255:0] testcases [7:0] = {
256'b0011000001001111110000001000000001100000000000011100001000000000000000001110000100000000000000000000000000000000000000000000010000110010000000010000000000000001000000011001100000000000000000000000110000010000000000000001111001000000000010010000111100000000, 256'b0110000111001001111011101000101000010010000011110010110010100100101011111011000100110110110011111100010110111000111011111110100111000010111100000000010111101011000001010101000111110011101010011001101000000100001100100010001101010110101110110100101110011000, 256'b0011000001001111110000001000000001100000000000011100001000000000000000001110000100000000000000000000000000000000000000000000010000110010000000010000000000000001000000011001100000000000000000000000110000010000000000000001111001000000000010010000111100000000, 256'b0110000111001001111011101000101000010010000011110010110010100100101011111011000100110110110011111100010110111000111011111110100111000010111100000000010111101011000001010101000111110011101010011001101000000100001100100010001101010110101110110100101110011000, 256'b0011111011000000010110110001111100000010111000011011111110100011000000011100000000010111101011000000000101000011110001101010001000101000000000000100000000000101010110101110110100000110001000010000011000000111011101000000000000000000001110000110000100000000, 256'b1111111111111111111111111111111111100011110111111111111111111111111111111111111111111111111111011111111111111111111111111101111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111111100111, 256'b001111101100000001011011000111110000001011100001101111111010001100000001110000000001011110101100000000010100001111000110101000100010100000000000010000000000010101011010111011010000011000100001000001100000011101110100000000000000000000101100011000010000000000000000, 256'b011111111111111111111111111111111110001111101111111111111111111111111111111111111111111111111101111111111111111111111111111011111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100101101111111111110011100000000
};
`endif
